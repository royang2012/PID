----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 11/12/2015 10:09:28 PM
-- Design Name: 
-- Module Name: log1215 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity log1215 is
    Port ( LOG_IN : in STD_LOGIC_VECTOR (11 downto 0);
           LOG_OUT : out STD_LOGIC_VECTOR (14 downto 0));
end log1215;

architecture Behavioral of log1215 is

begin
with LOG_IN select LOG_OUT <=
"000000000000000" when"000000000000",
"000000000000000" when"000000000001",
"000101010101011" when"000000000010",
"001000011101000" when"000000000011",
"001010101010101" when"000000000100",
"001100011000100" when"000000000101",
"001101110010011" when"000000000110",
"001110111110010" when"000000000111",
"010000000000000" when"000000001000",
"010000111010000" when"000000001001",
"010001101101111" when"000000001010",
"010010011100111" when"000000001011",
"010011000111101" when"000000001100",
"010011101111001" when"000000001101",
"010100010011101" when"000000001110",
"010100110101100" when"000000001111",
"010101010101011" when"000000010000",
"010101110011001" when"000000010001",
"010110001111011" when"000000010010",
"010110101010000" when"000000010011",
"010111000011010" when"000000010100",
"010111011011010" when"000000010101",
"010111110010001" when"000000010110",
"011000001000000" when"000000010111",
"011000011101000" when"000000011000",
"011000110001001" when"000000011001",
"011001000100011" when"000000011010",
"011001010111000" when"000000011011",
"011001101000111" when"000000011100",
"011001111010010" when"000000011101",
"011010001010111" when"000000011110",
"011010011011000" when"000000011111",
"011010101010101" when"000000100000",
"011010111001111" when"000000100001",
"011011001000100" when"000000100010",
"011011010110110" when"000000100011",
"011011100100101" when"000000100100",
"011011110010001" when"000000100101",
"011011111111010" when"000000100110",
"011100001100001" when"000000100111",
"011100011000100" when"000000101000",
"011100100100110" when"000000101001",
"011100110000101" when"000000101010",
"011100111100001" when"000000101011",
"011101000111100" when"000000101100",
"011101010010100" when"000000101101",
"011101011101011" when"000000101110",
"011101101000000" when"000000101111",
"011101110010011" when"000000110000",
"011101111100100" when"000000110001",
"011110000110011" when"000000110010",
"011110010000001" when"000000110011",
"011110011001110" when"000000110100",
"011110100011001" when"000000110101",
"011110101100011" when"000000110110",
"011110110101011" when"000000110111",
"011110111110010" when"000000111000",
"011111000111000" when"000000111001",
"011111001111100" when"000000111010",
"011111011000000" when"000000111011",
"011111100000010" when"000000111100",
"011111101000011" when"000000111101",
"011111110000011" when"000000111110",
"011111111000010" when"000000111111",
"100000000000000" when"000001000000",
"100000000111101" when"000001000001",
"100000001111001" when"000001000010",
"100000010110100" when"000001000011",
"100000011101111" when"000001000100",
"100000100101000" when"000001000101",
"100000101100001" when"000001000110",
"100000110011001" when"000001000111",
"100000111010000" when"000001001000",
"100001000000110" when"000001001001",
"100001000111100" when"000001001010",
"100001001110001" when"000001001011",
"100001010100101" when"000001001100",
"100001011011000" when"000001001101",
"100001100001011" when"000001001110",
"100001100111110" when"000001001111",
"100001101101111" when"000001010000",
"100001110100000" when"000001010001",
"100001111010000" when"000001010010",
"100010000000000" when"000001010011",
"100010000101111" when"000001010100",
"100010001011110" when"000001010101",
"100010010001100" when"000001010110",
"100010010111010" when"000001010111",
"100010011100111" when"000001011000",
"100010100010011" when"000001011001",
"100010100111111" when"000001011010",
"100010101101011" when"000001011011",
"100010110010110" when"000001011100",
"100010111000000" when"000001011101",
"100010111101010" when"000001011110",
"100011000010100" when"000001011111",
"100011000111101" when"000001100000",
"100011001100110" when"000001100001",
"100011010001111" when"000001100010",
"100011010110111" when"000001100011",
"100011011011110" when"000001100100",
"100011100000101" when"000001100101",
"100011100101100" when"000001100110",
"100011101010011" when"000001100111",
"100011101111001" when"000001101000",
"100011110011110" when"000001101001",
"100011111000100" when"000001101010",
"100011111101001" when"000001101011",
"100100000001101" when"000001101100",
"100100000110010" when"000001101101",
"100100001010110" when"000001101110",
"100100001111001" when"000001101111",
"100100010011101" when"000001110000",
"100100011000000" when"000001110001",
"100100011100010" when"000001110010",
"100100100000101" when"000001110011",
"100100100100111" when"000001110100",
"100100101001001" when"000001110101",
"100100101101010" when"000001110110",
"100100110001011" when"000001110111",
"100100110101100" when"000001111000",
"100100111001101" when"000001111001",
"100100111101110" when"000001111010",
"100101000001110" when"000001111011",
"100101000101110" when"000001111100",
"100101001001101" when"000001111101",
"100101001101101" when"000001111110",
"100101010001100" when"000001111111",
"100101010101011" when"000010000000",
"100101011001001" when"000010000001",
"100101011101000" when"000010000010",
"100101100000110" when"000010000011",
"100101100100100" when"000010000100",
"100101101000010" when"000010000101",
"100101101011111" when"000010000110",
"100101101111100" when"000010000111",
"100101110011001" when"000010001000",
"100101110110110" when"000010001001",
"100101111010011" when"000010001010",
"100101111101111" when"000010001011",
"100110000001100" when"000010001100",
"100110000101000" when"000010001101",
"100110001000100" when"000010001110",
"100110001011111" when"000010001111",
"100110001111011" when"000010010000",
"100110010010110" when"000010010001",
"100110010110001" when"000010010010",
"100110011001100" when"000010010011",
"100110011100111" when"000010010100",
"100110100000001" when"000010010101",
"100110100011011" when"000010010110",
"100110100110110" when"000010010111",
"100110101010000" when"000010011000",
"100110101101001" when"000010011001",
"100110110000011" when"000010011010",
"100110110011101" when"000010011011",
"100110110110110" when"000010011100",
"100110111001111" when"000010011101",
"100110111101000" when"000010011110",
"100111000000001" when"000010011111",
"100111000011010" when"000010100000",
"100111000110010" when"000010100001",
"100111001001011" when"000010100010",
"100111001100011" when"000010100011",
"100111001111011" when"000010100100",
"100111010010011" when"000010100101",
"100111010101011" when"000010100110",
"100111011000010" when"000010100111",
"100111011011010" when"000010101000",
"100111011110001" when"000010101001",
"100111100001001" when"000010101010",
"100111100100000" when"000010101011",
"100111100110111" when"000010101100",
"100111101001101" when"000010101101",
"100111101100100" when"000010101110",
"100111101111011" when"000010101111",
"100111110010001" when"000010110000",
"100111110101000" when"000010110001",
"100111110111110" when"000010110010",
"100111111010100" when"000010110011",
"100111111101010" when"000010110100",
"101000000000000" when"000010110101",
"101000000010101" when"000010110110",
"101000000101011" when"000010110111",
"101000001000000" when"000010111000",
"101000001010110" when"000010111001",
"101000001101011" when"000010111010",
"101000010000000" when"000010111011",
"101000010010101" when"000010111100",
"101000010101010" when"000010111101",
"101000010111111" when"000010111110",
"101000011010011" when"000010111111",
"101000011101000" when"000011000000",
"101000011111100" when"000011000001",
"101000100010001" when"000011000010",
"101000100100101" when"000011000011",
"101000100111001" when"000011000100",
"101000101001101" when"000011000101",
"101000101100001" when"000011000110",
"101000101110101" when"000011000111",
"101000110001001" when"000011001000",
"101000110011100" when"000011001001",
"101000110110000" when"000011001010",
"101000111000011" when"000011001011",
"101000111010111" when"000011001100",
"101000111101010" when"000011001101",
"101000111111101" when"000011001110",
"101001000010000" when"000011001111",
"101001000100011" when"000011010000",
"101001000110110" when"000011010001",
"101001001001001" when"000011010010",
"101001001011100" when"000011010011",
"101001001101110" when"000011010100",
"101001010000001" when"000011010101",
"101001010010011" when"000011010110",
"101001010100110" when"000011010111",
"101001010111000" when"000011011000",
"101001011001010" when"000011011001",
"101001011011100" when"000011011010",
"101001011101110" when"000011011011",
"101001100000000" when"000011011100",
"101001100010010" when"000011011101",
"101001100100100" when"000011011110",
"101001100110110" when"000011011111",
"101001101000111" when"000011100000",
"101001101011001" when"000011100001",
"101001101101010" when"000011100010",
"101001101111100" when"000011100011",
"101001110001101" when"000011100100",
"101001110011110" when"000011100101",
"101001110101111" when"000011100110",
"101001111000000" when"000011100111",
"101001111010010" when"000011101000",
"101001111100010" when"000011101001",
"101001111110011" when"000011101010",
"101010000000100" when"000011101011",
"101010000010101" when"000011101100",
"101010000100110" when"000011101101",
"101010000110110" when"000011101110",
"101010001000111" when"000011101111",
"101010001010111" when"000011110000",
"101010001100111" when"000011110001",
"101010001111000" when"000011110010",
"101010010001000" when"000011110011",
"101010010011000" when"000011110100",
"101010010101000" when"000011110101",
"101010010111000" when"000011110110",
"101010011001000" when"000011110111",
"101010011011000" when"000011111000",
"101010011101000" when"000011111001",
"101010011111000" when"000011111010",
"101010100001000" when"000011111011",
"101010100010111" when"000011111100",
"101010100100111" when"000011111101",
"101010100110110" when"000011111110",
"101010101000110" when"000011111111",
"101010101010101" when"000100000000",
"101010101100101" when"000100000001",
"101010101110100" when"000100000010",
"101010110000011" when"000100000011",
"101010110010010" when"000100000100",
"101010110100010" when"000100000101",
"101010110110001" when"000100000110",
"101010111000000" when"000100000111",
"101010111001111" when"000100001000",
"101010111011101" when"000100001001",
"101010111101100" when"000100001010",
"101010111111011" when"000100001011",
"101011000001010" when"000100001100",
"101011000011000" when"000100001101",
"101011000100111" when"000100001110",
"101011000110110" when"000100001111",
"101011001000100" when"000100010000",
"101011001010011" when"000100010001",
"101011001100001" when"000100010010",
"101011001101111" when"000100010011",
"101011001111110" when"000100010100",
"101011010001100" when"000100010101",
"101011010011010" when"000100010110",
"101011010101000" when"000100010111",
"101011010110110" when"000100011000",
"101011011000100" when"000100011001",
"101011011010010" when"000100011010",
"101011011100000" when"000100011011",
"101011011101110" when"000100011100",
"101011011111100" when"000100011101",
"101011100001010" when"000100011110",
"101011100011000" when"000100011111",
"101011100100101" when"000100100000",
"101011100110011" when"000100100001",
"101011101000001" when"000100100010",
"101011101001110" when"000100100011",
"101011101011100" when"000100100100",
"101011101101001" when"000100100101",
"101011101110111" when"000100100110",
"101011110000100" when"000100100111",
"101011110010001" when"000100101000",
"101011110011111" when"000100101001",
"101011110101100" when"000100101010",
"101011110111001" when"000100101011",
"101011111000110" when"000100101100",
"101011111010011" when"000100101101",
"101011111100000" when"000100101110",
"101011111101101" when"000100101111",
"101011111111010" when"000100110000",
"101100000000111" when"000100110001",
"101100000010100" when"000100110010",
"101100000100001" when"000100110011",
"101100000101110" when"000100110100",
"101100000111011" when"000100110101",
"101100001000111" when"000100110110",
"101100001010100" when"000100110111",
"101100001100001" when"000100111000",
"101100001101101" when"000100111001",
"101100001111010" when"000100111010",
"101100010000110" when"000100111011",
"101100010010011" when"000100111100",
"101100010011111" when"000100111101",
"101100010101100" when"000100111110",
"101100010111000" when"000100111111",
"101100011000100" when"000101000000",
"101100011010001" when"000101000001",
"101100011011101" when"000101000010",
"101100011101001" when"000101000011",
"101100011110101" when"000101000100",
"101100100000001" when"000101000101",
"101100100001110" when"000101000110",
"101100100011010" when"000101000111",
"101100100100110" when"000101001000",
"101100100110010" when"000101001001",
"101100100111110" when"000101001010",
"101100101001010" when"000101001011",
"101100101010101" when"000101001100",
"101100101100001" when"000101001101",
"101100101101101" when"000101001110",
"101100101111001" when"000101001111",
"101100110000101" when"000101010000",
"101100110010000" when"000101010001",
"101100110011100" when"000101010010",
"101100110101000" when"000101010011",
"101100110110011" when"000101010100",
"101100110111111" when"000101010101",
"101100111001010" when"000101010110",
"101100111010110" when"000101010111",
"101100111100001" when"000101011000",
"101100111101101" when"000101011001",
"101100111111000" when"000101011010",
"101101000000100" when"000101011011",
"101101000001111" when"000101011100",
"101101000011010" when"000101011101",
"101101000100101" when"000101011110",
"101101000110001" when"000101011111",
"101101000111100" when"000101100000",
"101101001000111" when"000101100001",
"101101001010010" when"000101100010",
"101101001011101" when"000101100011",
"101101001101000" when"000101100100",
"101101001110011" when"000101100101",
"101101001111110" when"000101100110",
"101101010001001" when"000101100111",
"101101010010100" when"000101101000",
"101101010011111" when"000101101001",
"101101010101010" when"000101101010",
"101101010110101" when"000101101011",
"101101011000000" when"000101101100",
"101101011001011" when"000101101101",
"101101011010110" when"000101101110",
"101101011100000" when"000101101111",
"101101011101011" when"000101110000",
"101101011110110" when"000101110001",
"101101100000000" when"000101110010",
"101101100001011" when"000101110011",
"101101100010110" when"000101110100",
"101101100100000" when"000101110101",
"101101100101011" when"000101110110",
"101101100110101" when"000101110111",
"101101101000000" when"000101111000",
"101101101001010" when"000101111001",
"101101101010101" when"000101111010",
"101101101011111" when"000101111011",
"101101101101001" when"000101111100",
"101101101110100" when"000101111101",
"101101101111110" when"000101111110",
"101101110001000" when"000101111111",
"101101110010011" when"000110000000",
"101101110011101" when"000110000001",
"101101110100111" when"000110000010",
"101101110110001" when"000110000011",
"101101110111011" when"000110000100",
"101101111000110" when"000110000101",
"101101111010000" when"000110000110",
"101101111011010" when"000110000111",
"101101111100100" when"000110001000",
"101101111101110" when"000110001001",
"101101111111000" when"000110001010",
"101110000000010" when"000110001011",
"101110000001100" when"000110001100",
"101110000010110" when"000110001101",
"101110000100000" when"000110001110",
"101110000101010" when"000110001111",
"101110000110011" when"000110010000",
"101110000111101" when"000110010001",
"101110001000111" when"000110010010",
"101110001010001" when"000110010011",
"101110001011011" when"000110010100",
"101110001100100" when"000110010101",
"101110001101110" when"000110010110",
"101110001111000" when"000110010111",
"101110010000001" when"000110011000",
"101110010001011" when"000110011001",
"101110010010101" when"000110011010",
"101110010011110" when"000110011011",
"101110010101000" when"000110011100",
"101110010110001" when"000110011101",
"101110010111011" when"000110011110",
"101110011000100" when"000110011111",
"101110011001110" when"000110100000",
"101110011010111" when"000110100001",
"101110011100001" when"000110100010",
"101110011101010" when"000110100011",
"101110011110100" when"000110100100",
"101110011111101" when"000110100101",
"101110100000110" when"000110100110",
"101110100010000" when"000110100111",
"101110100011001" when"000110101000",
"101110100100010" when"000110101001",
"101110100101100" when"000110101010",
"101110100110101" when"000110101011",
"101110100111110" when"000110101100",
"101110101000111" when"000110101101",
"101110101010000" when"000110101110",
"101110101011010" when"000110101111",
"101110101100011" when"000110110000",
"101110101101100" when"000110110001",
"101110101110101" when"000110110010",
"101110101111110" when"000110110011",
"101110110000111" when"000110110100",
"101110110010000" when"000110110101",
"101110110011001" when"000110110110",
"101110110100010" when"000110110111",
"101110110101011" when"000110111000",
"101110110110100" when"000110111001",
"101110110111101" when"000110111010",
"101110111000110" when"000110111011",
"101110111001111" when"000110111100",
"101110111010111" when"000110111101",
"101110111100000" when"000110111110",
"101110111101001" when"000110111111",
"101110111110010" when"000111000000",
"101110111111011" when"000111000001",
"101111000000011" when"000111000010",
"101111000001100" when"000111000011",
"101111000010101" when"000111000100",
"101111000011110" when"000111000101",
"101111000100110" when"000111000110",
"101111000101111" when"000111000111",
"101111000111000" when"000111001000",
"101111001000000" when"000111001001",
"101111001001001" when"000111001010",
"101111001010001" when"000111001011",
"101111001011010" when"000111001100",
"101111001100011" when"000111001101",
"101111001101011" when"000111001110",
"101111001110100" when"000111001111",
"101111001111100" when"000111010000",
"101111010000101" when"000111010001",
"101111010001101" when"000111010010",
"101111010010110" when"000111010011",
"101111010011110" when"000111010100",
"101111010100110" when"000111010101",
"101111010101111" when"000111010110",
"101111010110111" when"000111010111",
"101111011000000" when"000111011000",
"101111011001000" when"000111011001",
"101111011010000" when"000111011010",
"101111011011000" when"000111011011",
"101111011100001" when"000111011100",
"101111011101001" when"000111011101",
"101111011110001" when"000111011110",
"101111011111010" when"000111011111",
"101111100000010" when"000111100000",
"101111100001010" when"000111100001",
"101111100010010" when"000111100010",
"101111100011010" when"000111100011",
"101111100100010" when"000111100100",
"101111100101011" when"000111100101",
"101111100110011" when"000111100110",
"101111100111011" when"000111100111",
"101111101000011" when"000111101000",
"101111101001011" when"000111101001",
"101111101010011" when"000111101010",
"101111101011011" when"000111101011",
"101111101100011" when"000111101100",
"101111101101011" when"000111101101",
"101111101110011" when"000111101110",
"101111101111011" when"000111101111",
"101111110000011" when"000111110000",
"101111110001011" when"000111110001",
"101111110010011" when"000111110010",
"101111110011011" when"000111110011",
"101111110100011" when"000111110100",
"101111110101010" when"000111110101",
"101111110110010" when"000111110110",
"101111110111010" when"000111110111",
"101111111000010" when"000111111000",
"101111111001010" when"000111111001",
"101111111010010" when"000111111010",
"101111111011001" when"000111111011",
"101111111100001" when"000111111100",
"101111111101001" when"000111111101",
"101111111110001" when"000111111110",
"101111111111000" when"000111111111",
"110000000000000" when"001000000000",
"110000000001000" when"001000000001",
"110000000001111" when"001000000010",
"110000000010111" when"001000000011",
"110000000011111" when"001000000100",
"110000000100110" when"001000000101",
"110000000101110" when"001000000110",
"110000000110101" when"001000000111",
"110000000111101" when"001000001000",
"110000001000101" when"001000001001",
"110000001001100" when"001000001010",
"110000001010100" when"001000001011",
"110000001011011" when"001000001100",
"110000001100011" when"001000001101",
"110000001101010" when"001000001110",
"110000001110010" when"001000001111",
"110000001111001" when"001000010000",
"110000010000001" when"001000010001",
"110000010001000" when"001000010010",
"110000010010000" when"001000010011",
"110000010010111" when"001000010100",
"110000010011110" when"001000010101",
"110000010100110" when"001000010110",
"110000010101101" when"001000010111",
"110000010110100" when"001000011000",
"110000010111100" when"001000011001",
"110000011000011" when"001000011010",
"110000011001010" when"001000011011",
"110000011010010" when"001000011100",
"110000011011001" when"001000011101",
"110000011100000" when"001000011110",
"110000011101000" when"001000011111",
"110000011101111" when"001000100000",
"110000011110110" when"001000100001",
"110000011111101" when"001000100010",
"110000100000100" when"001000100011",
"110000100001100" when"001000100100",
"110000100010011" when"001000100101",
"110000100011010" when"001000100110",
"110000100100001" when"001000100111",
"110000100101000" when"001000101000",
"110000100101111" when"001000101001",
"110000100110111" when"001000101010",
"110000100111110" when"001000101011",
"110000101000101" when"001000101100",
"110000101001100" when"001000101101",
"110000101010011" when"001000101110",
"110000101011010" when"001000101111",
"110000101100001" when"001000110000",
"110000101101000" when"001000110001",
"110000101101111" when"001000110010",
"110000101110110" when"001000110011",
"110000101111101" when"001000110100",
"110000110000100" when"001000110101",
"110000110001011" when"001000110110",
"110000110010010" when"001000110111",
"110000110011001" when"001000111000",
"110000110100000" when"001000111001",
"110000110100111" when"001000111010",
"110000110101110" when"001000111011",
"110000110110101" when"001000111100",
"110000110111011" when"001000111101",
"110000111000010" when"001000111110",
"110000111001001" when"001000111111",
"110000111010000" when"001001000000",
"110000111010111" when"001001000001",
"110000111011110" when"001001000010",
"110000111100100" when"001001000011",
"110000111101011" when"001001000100",
"110000111110010" when"001001000101",
"110000111111001" when"001001000110",
"110001000000000" when"001001000111",
"110001000000110" when"001001001000",
"110001000001101" when"001001001001",
"110001000010100" when"001001001010",
"110001000011011" when"001001001011",
"110001000100001" when"001001001100",
"110001000101000" when"001001001101",
"110001000101111" when"001001001110",
"110001000110101" when"001001001111",
"110001000111100" when"001001010000",
"110001001000011" when"001001010001",
"110001001001001" when"001001010010",
"110001001010000" when"001001010011",
"110001001010110" when"001001010100",
"110001001011101" when"001001010101",
"110001001100100" when"001001010110",
"110001001101010" when"001001010111",
"110001001110001" when"001001011000",
"110001001110111" when"001001011001",
"110001001111110" when"001001011010",
"110001010000100" when"001001011011",
"110001010001011" when"001001011100",
"110001010010001" when"001001011101",
"110001010011000" when"001001011110",
"110001010011110" when"001001011111",
"110001010100101" when"001001100000",
"110001010101011" when"001001100001",
"110001010110010" when"001001100010",
"110001010111000" when"001001100011",
"110001010111111" when"001001100100",
"110001011000101" when"001001100101",
"110001011001100" when"001001100110",
"110001011010010" when"001001100111",
"110001011011000" when"001001101000",
"110001011011111" when"001001101001",
"110001011100101" when"001001101010",
"110001011101100" when"001001101011",
"110001011110010" when"001001101100",
"110001011111000" when"001001101101",
"110001011111111" when"001001101110",
"110001100000101" when"001001101111",
"110001100001011" when"001001110000",
"110001100010010" when"001001110001",
"110001100011000" when"001001110010",
"110001100011110" when"001001110011",
"110001100100100" when"001001110100",
"110001100101011" when"001001110101",
"110001100110001" when"001001110110",
"110001100110111" when"001001110111",
"110001100111101" when"001001111000",
"110001101000100" when"001001111001",
"110001101001010" when"001001111010",
"110001101010000" when"001001111011",
"110001101010110" when"001001111100",
"110001101011101" when"001001111101",
"110001101100011" when"001001111110",
"110001101101001" when"001001111111",
"110001101101111" when"001010000000",
"110001101110101" when"001010000001",
"110001101111011" when"001010000010",
"110001110000001" when"001010000011",
"110001110001000" when"001010000100",
"110001110001110" when"001010000101",
"110001110010100" when"001010000110",
"110001110011010" when"001010000111",
"110001110100000" when"001010001000",
"110001110100110" when"001010001001",
"110001110101100" when"001010001010",
"110001110110010" when"001010001011",
"110001110111000" when"001010001100",
"110001110111110" when"001010001101",
"110001111000100" when"001010001110",
"110001111001010" when"001010001111",
"110001111010000" when"001010010000",
"110001111010110" when"001010010001",
"110001111011100" when"001010010010",
"110001111100010" when"001010010011",
"110001111101000" when"001010010100",
"110001111101110" when"001010010101",
"110001111110100" when"001010010110",
"110001111111010" when"001010010111",
"110010000000000" when"001010011000",
"110010000000110" when"001010011001",
"110010000001100" when"001010011010",
"110010000010010" when"001010011011",
"110010000011000" when"001010011100",
"110010000011110" when"001010011101",
"110010000100100" when"001010011110",
"110010000101001" when"001010011111",
"110010000101111" when"001010100000",
"110010000110101" when"001010100001",
"110010000111011" when"001010100010",
"110010001000001" when"001010100011",
"110010001000111" when"001010100100",
"110010001001100" when"001010100101",
"110010001010010" when"001010100110",
"110010001011000" when"001010100111",
"110010001011110" when"001010101000",
"110010001100100" when"001010101001",
"110010001101001" when"001010101010",
"110010001101111" when"001010101011",
"110010001110101" when"001010101100",
"110010001111011" when"001010101101",
"110010010000000" when"001010101110",
"110010010000110" when"001010101111",
"110010010001100" when"001010110000",
"110010010010010" when"001010110001",
"110010010010111" when"001010110010",
"110010010011101" when"001010110011",
"110010010100011" when"001010110100",
"110010010101000" when"001010110101",
"110010010101110" when"001010110110",
"110010010110100" when"001010110111",
"110010010111010" when"001010111000",
"110010010111111" when"001010111001",
"110010011000101" when"001010111010",
"110010011001010" when"001010111011",
"110010011010000" when"001010111100",
"110010011010110" when"001010111101",
"110010011011011" when"001010111110",
"110010011100001" when"001010111111",
"110010011100111" when"001011000000",
"110010011101100" when"001011000001",
"110010011110010" when"001011000010",
"110010011110111" when"001011000011",
"110010011111101" when"001011000100",
"110010100000010" when"001011000101",
"110010100001000" when"001011000110",
"110010100001110" when"001011000111",
"110010100010011" when"001011001000",
"110010100011001" when"001011001001",
"110010100011110" when"001011001010",
"110010100100100" when"001011001011",
"110010100101001" when"001011001100",
"110010100101111" when"001011001101",
"110010100110100" when"001011001110",
"110010100111010" when"001011001111",
"110010100111111" when"001011010000",
"110010101000101" when"001011010001",
"110010101001010" when"001011010010",
"110010101001111" when"001011010011",
"110010101010101" when"001011010100",
"110010101011010" when"001011010101",
"110010101100000" when"001011010110",
"110010101100101" when"001011010111",
"110010101101011" when"001011011000",
"110010101110000" when"001011011001",
"110010101110101" when"001011011010",
"110010101111011" when"001011011011",
"110010110000000" when"001011011100",
"110010110000110" when"001011011101",
"110010110001011" when"001011011110",
"110010110010000" when"001011011111",
"110010110010110" when"001011100000",
"110010110011011" when"001011100001",
"110010110100000" when"001011100010",
"110010110100110" when"001011100011",
"110010110101011" when"001011100100",
"110010110110000" when"001011100101",
"110010110110110" when"001011100110",
"110010110111011" when"001011100111",
"110010111000000" when"001011101000",
"110010111000110" when"001011101001",
"110010111001011" when"001011101010",
"110010111010000" when"001011101011",
"110010111010101" when"001011101100",
"110010111011011" when"001011101101",
"110010111100000" when"001011101110",
"110010111100101" when"001011101111",
"110010111101010" when"001011110000",
"110010111110000" when"001011110001",
"110010111110101" when"001011110010",
"110010111111010" when"001011110011",
"110010111111111" when"001011110100",
"110011000000100" when"001011110101",
"110011000001010" when"001011110110",
"110011000001111" when"001011110111",
"110011000010100" when"001011111000",
"110011000011001" when"001011111001",
"110011000011110" when"001011111010",
"110011000100100" when"001011111011",
"110011000101001" when"001011111100",
"110011000101110" when"001011111101",
"110011000110011" when"001011111110",
"110011000111000" when"001011111111",
"110011000111101" when"001100000000",
"110011001000010" when"001100000001",
"110011001001000" when"001100000010",
"110011001001101" when"001100000011",
"110011001010010" when"001100000100",
"110011001010111" when"001100000101",
"110011001011100" when"001100000110",
"110011001100001" when"001100000111",
"110011001100110" when"001100001000",
"110011001101011" when"001100001001",
"110011001110000" when"001100001010",
"110011001110101" when"001100001011",
"110011001111010" when"001100001100",
"110011001111111" when"001100001101",
"110011010000100" when"001100001110",
"110011010001010" when"001100001111",
"110011010001111" when"001100010000",
"110011010010100" when"001100010001",
"110011010011001" when"001100010010",
"110011010011110" when"001100010011",
"110011010100011" when"001100010100",
"110011010101000" when"001100010101",
"110011010101101" when"001100010110",
"110011010110010" when"001100010111",
"110011010110111" when"001100011000",
"110011010111100" when"001100011001",
"110011011000000" when"001100011010",
"110011011000101" when"001100011011",
"110011011001010" when"001100011100",
"110011011001111" when"001100011101",
"110011011010100" when"001100011110",
"110011011011001" when"001100011111",
"110011011011110" when"001100100000",
"110011011100011" when"001100100001",
"110011011101000" when"001100100010",
"110011011101101" when"001100100011",
"110011011110010" when"001100100100",
"110011011110111" when"001100100101",
"110011011111100" when"001100100110",
"110011100000000" when"001100100111",
"110011100000101" when"001100101000",
"110011100001010" when"001100101001",
"110011100001111" when"001100101010",
"110011100010100" when"001100101011",
"110011100011001" when"001100101100",
"110011100011110" when"001100101101",
"110011100100010" when"001100101110",
"110011100100111" when"001100101111",
"110011100101100" when"001100110000",
"110011100110001" when"001100110001",
"110011100110110" when"001100110010",
"110011100111011" when"001100110011",
"110011100111111" when"001100110100",
"110011101000100" when"001100110101",
"110011101001001" when"001100110110",
"110011101001110" when"001100110111",
"110011101010011" when"001100111000",
"110011101010111" when"001100111001",
"110011101011100" when"001100111010",
"110011101100001" when"001100111011",
"110011101100110" when"001100111100",
"110011101101010" when"001100111101",
"110011101101111" when"001100111110",
"110011101110100" when"001100111111",
"110011101111001" when"001101000000",
"110011101111101" when"001101000001",
"110011110000010" when"001101000010",
"110011110000111" when"001101000011",
"110011110001100" when"001101000100",
"110011110010000" when"001101000101",
"110011110010101" when"001101000110",
"110011110011010" when"001101000111",
"110011110011110" when"001101001000",
"110011110100011" when"001101001001",
"110011110101000" when"001101001010",
"110011110101100" when"001101001011",
"110011110110001" when"001101001100",
"110011110110110" when"001101001101",
"110011110111010" when"001101001110",
"110011110111111" when"001101001111",
"110011111000100" when"001101010000",
"110011111001000" when"001101010001",
"110011111001101" when"001101010010",
"110011111010010" when"001101010011",
"110011111010110" when"001101010100",
"110011111011011" when"001101010101",
"110011111011111" when"001101010110",
"110011111100100" when"001101010111",
"110011111101001" when"001101011000",
"110011111101101" when"001101011001",
"110011111110010" when"001101011010",
"110011111110110" when"001101011011",
"110011111111011" when"001101011100",
"110100000000000" when"001101011101",
"110100000000100" when"001101011110",
"110100000001001" when"001101011111",
"110100000001101" when"001101100000",
"110100000010010" when"001101100001",
"110100000010110" when"001101100010",
"110100000011011" when"001101100011",
"110100000100000" when"001101100100",
"110100000100100" when"001101100101",
"110100000101001" when"001101100110",
"110100000101101" when"001101100111",
"110100000110010" when"001101101000",
"110100000110110" when"001101101001",
"110100000111011" when"001101101010",
"110100000111111" when"001101101011",
"110100001000100" when"001101101100",
"110100001001000" when"001101101101",
"110100001001101" when"001101101110",
"110100001010001" when"001101101111",
"110100001010110" when"001101110000",
"110100001011010" when"001101110001",
"110100001011111" when"001101110010",
"110100001100011" when"001101110011",
"110100001100111" when"001101110100",
"110100001101100" when"001101110101",
"110100001110000" when"001101110110",
"110100001110101" when"001101110111",
"110100001111001" when"001101111000",
"110100001111110" when"001101111001",
"110100010000010" when"001101111010",
"110100010000111" when"001101111011",
"110100010001011" when"001101111100",
"110100010001111" when"001101111101",
"110100010010100" when"001101111110",
"110100010011000" when"001101111111",
"110100010011101" when"001110000000",
"110100010100001" when"001110000001",
"110100010100101" when"001110000010",
"110100010101010" when"001110000011",
"110100010101110" when"001110000100",
"110100010110011" when"001110000101",
"110100010110111" when"001110000110",
"110100010111011" when"001110000111",
"110100011000000" when"001110001000",
"110100011000100" when"001110001001",
"110100011001000" when"001110001010",
"110100011001101" when"001110001011",
"110100011010001" when"001110001100",
"110100011010101" when"001110001101",
"110100011011010" when"001110001110",
"110100011011110" when"001110001111",
"110100011100010" when"001110010000",
"110100011100111" when"001110010001",
"110100011101011" when"001110010010",
"110100011101111" when"001110010011",
"110100011110100" when"001110010100",
"110100011111000" when"001110010101",
"110100011111100" when"001110010110",
"110100100000000" when"001110010111",
"110100100000101" when"001110011000",
"110100100001001" when"001110011001",
"110100100001101" when"001110011010",
"110100100010010" when"001110011011",
"110100100010110" when"001110011100",
"110100100011010" when"001110011101",
"110100100011110" when"001110011110",
"110100100100011" when"001110011111",
"110100100100111" when"001110100000",
"110100100101011" when"001110100001",
"110100100101111" when"001110100010",
"110100100110100" when"001110100011",
"110100100111000" when"001110100100",
"110100100111100" when"001110100101",
"110100101000000" when"001110100110",
"110100101000100" when"001110100111",
"110100101001001" when"001110101000",
"110100101001101" when"001110101001",
"110100101010001" when"001110101010",
"110100101010101" when"001110101011",
"110100101011001" when"001110101100",
"110100101011110" when"001110101101",
"110100101100010" when"001110101110",
"110100101100110" when"001110101111",
"110100101101010" when"001110110000",
"110100101101110" when"001110110001",
"110100101110011" when"001110110010",
"110100101110111" when"001110110011",
"110100101111011" when"001110110100",
"110100101111111" when"001110110101",
"110100110000011" when"001110110110",
"110100110000111" when"001110110111",
"110100110001011" when"001110111000",
"110100110010000" when"001110111001",
"110100110010100" when"001110111010",
"110100110011000" when"001110111011",
"110100110011100" when"001110111100",
"110100110100000" when"001110111101",
"110100110100100" when"001110111110",
"110100110101000" when"001110111111",
"110100110101100" when"001111000000",
"110100110110000" when"001111000001",
"110100110110101" when"001111000010",
"110100110111001" when"001111000011",
"110100110111101" when"001111000100",
"110100111000001" when"001111000101",
"110100111000101" when"001111000110",
"110100111001001" when"001111000111",
"110100111001101" when"001111001000",
"110100111010001" when"001111001001",
"110100111010101" when"001111001010",
"110100111011001" when"001111001011",
"110100111011101" when"001111001100",
"110100111100001" when"001111001101",
"110100111100101" when"001111001110",
"110100111101001" when"001111001111",
"110100111101110" when"001111010000",
"110100111110010" when"001111010001",
"110100111110110" when"001111010010",
"110100111111010" when"001111010011",
"110100111111110" when"001111010100",
"110101000000010" when"001111010101",
"110101000000110" when"001111010110",
"110101000001010" when"001111010111",
"110101000001110" when"001111011000",
"110101000010010" when"001111011001",
"110101000010110" when"001111011010",
"110101000011010" when"001111011011",
"110101000011110" when"001111011100",
"110101000100010" when"001111011101",
"110101000100110" when"001111011110",
"110101000101010" when"001111011111",
"110101000101110" when"001111100000",
"110101000110010" when"001111100001",
"110101000110101" when"001111100010",
"110101000111001" when"001111100011",
"110101000111101" when"001111100100",
"110101001000001" when"001111100101",
"110101001000101" when"001111100110",
"110101001001001" when"001111100111",
"110101001001101" when"001111101000",
"110101001010001" when"001111101001",
"110101001010101" when"001111101010",
"110101001011001" when"001111101011",
"110101001011101" when"001111101100",
"110101001100001" when"001111101101",
"110101001100101" when"001111101110",
"110101001101001" when"001111101111",
"110101001101101" when"001111110000",
"110101001110001" when"001111110001",
"110101001110100" when"001111110010",
"110101001111000" when"001111110011",
"110101001111100" when"001111110100",
"110101010000000" when"001111110101",
"110101010000100" when"001111110110",
"110101010001000" when"001111110111",
"110101010001100" when"001111111000",
"110101010010000" when"001111111001",
"110101010010011" when"001111111010",
"110101010010111" when"001111111011",
"110101010011011" when"001111111100",
"110101010011111" when"001111111101",
"110101010100011" when"001111111110",
"110101010100111" when"001111111111",
"110101010101011" when"010000000000",
"110101010101110" when"010000000001",
"110101010110010" when"010000000010",
"110101010110110" when"010000000011",
"110101010111010" when"010000000100",
"110101010111110" when"010000000101",
"110101011000010" when"010000000110",
"110101011000101" when"010000000111",
"110101011001001" when"010000001000",
"110101011001101" when"010000001001",
"110101011010001" when"010000001010",
"110101011010101" when"010000001011",
"110101011011001" when"010000001100",
"110101011011100" when"010000001101",
"110101011100000" when"010000001110",
"110101011100100" when"010000001111",
"110101011101000" when"010000010000",
"110101011101100" when"010000010001",
"110101011101111" when"010000010010",
"110101011110011" when"010000010011",
"110101011110111" when"010000010100",
"110101011111011" when"010000010101",
"110101011111110" when"010000010110",
"110101100000010" when"010000010111",
"110101100000110" when"010000011000",
"110101100001010" when"010000011001",
"110101100001101" when"010000011010",
"110101100010001" when"010000011011",
"110101100010101" when"010000011100",
"110101100011001" when"010000011101",
"110101100011100" when"010000011110",
"110101100100000" when"010000011111",
"110101100100100" when"010000100000",
"110101100101000" when"010000100001",
"110101100101011" when"010000100010",
"110101100101111" when"010000100011",
"110101100110011" when"010000100100",
"110101100110110" when"010000100101",
"110101100111010" when"010000100110",
"110101100111110" when"010000100111",
"110101101000010" when"010000101000",
"110101101000101" when"010000101001",
"110101101001001" when"010000101010",
"110101101001101" when"010000101011",
"110101101010000" when"010000101100",
"110101101010100" when"010000101101",
"110101101011000" when"010000101110",
"110101101011011" when"010000101111",
"110101101011111" when"010000110000",
"110101101100011" when"010000110001",
"110101101100110" when"010000110010",
"110101101101010" when"010000110011",
"110101101101110" when"010000110100",
"110101101110001" when"010000110101",
"110101101110101" when"010000110110",
"110101101111001" when"010000110111",
"110101101111100" when"010000111000",
"110101110000000" when"010000111001",
"110101110000100" when"010000111010",
"110101110000111" when"010000111011",
"110101110001011" when"010000111100",
"110101110001111" when"010000111101",
"110101110010010" when"010000111110",
"110101110010110" when"010000111111",
"110101110011001" when"010001000000",
"110101110011101" when"010001000001",
"110101110100001" when"010001000010",
"110101110100100" when"010001000011",
"110101110101000" when"010001000100",
"110101110101100" when"010001000101",
"110101110101111" when"010001000110",
"110101110110011" when"010001000111",
"110101110110110" when"010001001000",
"110101110111010" when"010001001001",
"110101110111110" when"010001001010",
"110101111000001" when"010001001011",
"110101111000101" when"010001001100",
"110101111001000" when"010001001101",
"110101111001100" when"010001001110",
"110101111001111" when"010001001111",
"110101111010011" when"010001010000",
"110101111010111" when"010001010001",
"110101111011010" when"010001010010",
"110101111011110" when"010001010011",
"110101111100001" when"010001010100",
"110101111100101" when"010001010101",
"110101111101000" when"010001010110",
"110101111101100" when"010001010111",
"110101111101111" when"010001011000",
"110101111110011" when"010001011001",
"110101111110111" when"010001011010",
"110101111111010" when"010001011011",
"110101111111110" when"010001011100",
"110110000000001" when"010001011101",
"110110000000101" when"010001011110",
"110110000001000" when"010001011111",
"110110000001100" when"010001100000",
"110110000001111" when"010001100001",
"110110000010011" when"010001100010",
"110110000010110" when"010001100011",
"110110000011010" when"010001100100",
"110110000011101" when"010001100101",
"110110000100001" when"010001100110",
"110110000100100" when"010001100111",
"110110000101000" when"010001101000",
"110110000101011" when"010001101001",
"110110000101111" when"010001101010",
"110110000110010" when"010001101011",
"110110000110110" when"010001101100",
"110110000111001" when"010001101101",
"110110000111101" when"010001101110",
"110110001000000" when"010001101111",
"110110001000100" when"010001110000",
"110110001000111" when"010001110001",
"110110001001010" when"010001110010",
"110110001001110" when"010001110011",
"110110001010001" when"010001110100",
"110110001010101" when"010001110101",
"110110001011000" when"010001110110",
"110110001011100" when"010001110111",
"110110001011111" when"010001111000",
"110110001100011" when"010001111001",
"110110001100110" when"010001111010",
"110110001101010" when"010001111011",
"110110001101101" when"010001111100",
"110110001110000" when"010001111101",
"110110001110100" when"010001111110",
"110110001110111" when"010001111111",
"110110001111011" when"010010000000",
"110110001111110" when"010010000001",
"110110010000001" when"010010000010",
"110110010000101" when"010010000011",
"110110010001000" when"010010000100",
"110110010001100" when"010010000101",
"110110010001111" when"010010000110",
"110110010010011" when"010010000111",
"110110010010110" when"010010001000",
"110110010011001" when"010010001001",
"110110010011101" when"010010001010",
"110110010100000" when"010010001011",
"110110010100011" when"010010001100",
"110110010100111" when"010010001101",
"110110010101010" when"010010001110",
"110110010101110" when"010010001111",
"110110010110001" when"010010010000",
"110110010110100" when"010010010001",
"110110010111000" when"010010010010",
"110110010111011" when"010010010011",
"110110010111110" when"010010010100",
"110110011000010" when"010010010101",
"110110011000101" when"010010010110",
"110110011001001" when"010010010111",
"110110011001100" when"010010011000",
"110110011001111" when"010010011001",
"110110011010011" when"010010011010",
"110110011010110" when"010010011011",
"110110011011001" when"010010011100",
"110110011011101" when"010010011101",
"110110011100000" when"010010011110",
"110110011100011" when"010010011111",
"110110011100111" when"010010100000",
"110110011101010" when"010010100001",
"110110011101101" when"010010100010",
"110110011110001" when"010010100011",
"110110011110100" when"010010100100",
"110110011110111" when"010010100101",
"110110011111010" when"010010100110",
"110110011111110" when"010010100111",
"110110100000001" when"010010101000",
"110110100000100" when"010010101001",
"110110100001000" when"010010101010",
"110110100001011" when"010010101011",
"110110100001110" when"010010101100",
"110110100010010" when"010010101101",
"110110100010101" when"010010101110",
"110110100011000" when"010010101111",
"110110100011011" when"010010110000",
"110110100011111" when"010010110001",
"110110100100010" when"010010110010",
"110110100100101" when"010010110011",
"110110100101001" when"010010110100",
"110110100101100" when"010010110101",
"110110100101111" when"010010110110",
"110110100110010" when"010010110111",
"110110100110110" when"010010111000",
"110110100111001" when"010010111001",
"110110100111100" when"010010111010",
"110110100111111" when"010010111011",
"110110101000011" when"010010111100",
"110110101000110" when"010010111101",
"110110101001001" when"010010111110",
"110110101001100" when"010010111111",
"110110101010000" when"010011000000",
"110110101010011" when"010011000001",
"110110101010110" when"010011000010",
"110110101011001" when"010011000011",
"110110101011101" when"010011000100",
"110110101100000" when"010011000101",
"110110101100011" when"010011000110",
"110110101100110" when"010011000111",
"110110101101001" when"010011001000",
"110110101101101" when"010011001001",
"110110101110000" when"010011001010",
"110110101110011" when"010011001011",
"110110101110110" when"010011001100",
"110110101111010" when"010011001101",
"110110101111101" when"010011001110",
"110110110000000" when"010011001111",
"110110110000011" when"010011010000",
"110110110000110" when"010011010001",
"110110110001010" when"010011010010",
"110110110001101" when"010011010011",
"110110110010000" when"010011010100",
"110110110010011" when"010011010101",
"110110110010110" when"010011010110",
"110110110011001" when"010011010111",
"110110110011101" when"010011011000",
"110110110100000" when"010011011001",
"110110110100011" when"010011011010",
"110110110100110" when"010011011011",
"110110110101001" when"010011011100",
"110110110101100" when"010011011101",
"110110110110000" when"010011011110",
"110110110110011" when"010011011111",
"110110110110110" when"010011100000",
"110110110111001" when"010011100001",
"110110110111100" when"010011100010",
"110110110111111" when"010011100011",
"110110111000011" when"010011100100",
"110110111000110" when"010011100101",
"110110111001001" when"010011100110",
"110110111001100" when"010011100111",
"110110111001111" when"010011101000",
"110110111010010" when"010011101001",
"110110111010101" when"010011101010",
"110110111011001" when"010011101011",
"110110111011100" when"010011101100",
"110110111011111" when"010011101101",
"110110111100010" when"010011101110",
"110110111100101" when"010011101111",
"110110111101000" when"010011110000",
"110110111101011" when"010011110001",
"110110111101110" when"010011110010",
"110110111110001" when"010011110011",
"110110111110101" when"010011110100",
"110110111111000" when"010011110101",
"110110111111011" when"010011110110",
"110110111111110" when"010011110111",
"110111000000001" when"010011111000",
"110111000000100" when"010011111001",
"110111000000111" when"010011111010",
"110111000001010" when"010011111011",
"110111000001101" when"010011111100",
"110111000010000" when"010011111101",
"110111000010100" when"010011111110",
"110111000010111" when"010011111111",
"110111000011010" when"010100000000",
"110111000011101" when"010100000001",
"110111000100000" when"010100000010",
"110111000100011" when"010100000011",
"110111000100110" when"010100000100",
"110111000101001" when"010100000101",
"110111000101100" when"010100000110",
"110111000101111" when"010100000111",
"110111000110010" when"010100001000",
"110111000110101" when"010100001001",
"110111000111000" when"010100001010",
"110111000111011" when"010100001011",
"110111000111110" when"010100001100",
"110111001000010" when"010100001101",
"110111001000101" when"010100001110",
"110111001001000" when"010100001111",
"110111001001011" when"010100010000",
"110111001001110" when"010100010001",
"110111001010001" when"010100010010",
"110111001010100" when"010100010011",
"110111001010111" when"010100010100",
"110111001011010" when"010100010101",
"110111001011101" when"010100010110",
"110111001100000" when"010100010111",
"110111001100011" when"010100011000",
"110111001100110" when"010100011001",
"110111001101001" when"010100011010",
"110111001101100" when"010100011011",
"110111001101111" when"010100011100",
"110111001110010" when"010100011101",
"110111001110101" when"010100011110",
"110111001111000" when"010100011111",
"110111001111011" when"010100100000",
"110111001111110" when"010100100001",
"110111010000001" when"010100100010",
"110111010000100" when"010100100011",
"110111010000111" when"010100100100",
"110111010001010" when"010100100101",
"110111010001101" when"010100100110",
"110111010010000" when"010100100111",
"110111010010011" when"010100101000",
"110111010010110" when"010100101001",
"110111010011001" when"010100101010",
"110111010011100" when"010100101011",
"110111010011111" when"010100101100",
"110111010100010" when"010100101101",
"110111010100101" when"010100101110",
"110111010101000" when"010100101111",
"110111010101011" when"010100110000",
"110111010101110" when"010100110001",
"110111010110001" when"010100110010",
"110111010110100" when"010100110011",
"110111010110111" when"010100110100",
"110111010111010" when"010100110101",
"110111010111101" when"010100110110",
"110111010111111" when"010100110111",
"110111011000010" when"010100111000",
"110111011000101" when"010100111001",
"110111011001000" when"010100111010",
"110111011001011" when"010100111011",
"110111011001110" when"010100111100",
"110111011010001" when"010100111101",
"110111011010100" when"010100111110",
"110111011010111" when"010100111111",
"110111011011010" when"010101000000",
"110111011011101" when"010101000001",
"110111011100000" when"010101000010",
"110111011100011" when"010101000011",
"110111011100110" when"010101000100",
"110111011101001" when"010101000101",
"110111011101011" when"010101000110",
"110111011101110" when"010101000111",
"110111011110001" when"010101001000",
"110111011110100" when"010101001001",
"110111011110111" when"010101001010",
"110111011111010" when"010101001011",
"110111011111101" when"010101001100",
"110111100000000" when"010101001101",
"110111100000011" when"010101001110",
"110111100000110" when"010101001111",
"110111100001001" when"010101010000",
"110111100001011" when"010101010001",
"110111100001110" when"010101010010",
"110111100010001" when"010101010011",
"110111100010100" when"010101010100",
"110111100010111" when"010101010101",
"110111100011010" when"010101010110",
"110111100011101" when"010101010111",
"110111100100000" when"010101011000",
"110111100100011" when"010101011001",
"110111100100101" when"010101011010",
"110111100101000" when"010101011011",
"110111100101011" when"010101011100",
"110111100101110" when"010101011101",
"110111100110001" when"010101011110",
"110111100110100" when"010101011111",
"110111100110111" when"010101100000",
"110111100111001" when"010101100001",
"110111100111100" when"010101100010",
"110111100111111" when"010101100011",
"110111101000010" when"010101100100",
"110111101000101" when"010101100101",
"110111101001000" when"010101100110",
"110111101001011" when"010101100111",
"110111101001101" when"010101101000",
"110111101010000" when"010101101001",
"110111101010011" when"010101101010",
"110111101010110" when"010101101011",
"110111101011001" when"010101101100",
"110111101011100" when"010101101101",
"110111101011111" when"010101101110",
"110111101100001" when"010101101111",
"110111101100100" when"010101110000",
"110111101100111" when"010101110001",
"110111101101010" when"010101110010",
"110111101101101" when"010101110011",
"110111101101111" when"010101110100",
"110111101110010" when"010101110101",
"110111101110101" when"010101110110",
"110111101111000" when"010101110111",
"110111101111011" when"010101111000",
"110111101111110" when"010101111001",
"110111110000000" when"010101111010",
"110111110000011" when"010101111011",
"110111110000110" when"010101111100",
"110111110001001" when"010101111101",
"110111110001100" when"010101111110",
"110111110001110" when"010101111111",
"110111110010001" when"010110000000",
"110111110010100" when"010110000001",
"110111110010111" when"010110000010",
"110111110011010" when"010110000011",
"110111110011100" when"010110000100",
"110111110011111" when"010110000101",
"110111110100010" when"010110000110",
"110111110100101" when"010110000111",
"110111110101000" when"010110001000",
"110111110101010" when"010110001001",
"110111110101101" when"010110001010",
"110111110110000" when"010110001011",
"110111110110011" when"010110001100",
"110111110110101" when"010110001101",
"110111110111000" when"010110001110",
"110111110111011" when"010110001111",
"110111110111110" when"010110010000",
"110111111000000" when"010110010001",
"110111111000011" when"010110010010",
"110111111000110" when"010110010011",
"110111111001001" when"010110010100",
"110111111001100" when"010110010101",
"110111111001110" when"010110010110",
"110111111010001" when"010110010111",
"110111111010100" when"010110011000",
"110111111010111" when"010110011001",
"110111111011001" when"010110011010",
"110111111011100" when"010110011011",
"110111111011111" when"010110011100",
"110111111100010" when"010110011101",
"110111111100100" when"010110011110",
"110111111100111" when"010110011111",
"110111111101010" when"010110100000",
"110111111101100" when"010110100001",
"110111111101111" when"010110100010",
"110111111110010" when"010110100011",
"110111111110101" when"010110100100",
"110111111110111" when"010110100101",
"110111111111010" when"010110100110",
"110111111111101" when"010110100111",
"111000000000000" when"010110101000",
"111000000000010" when"010110101001",
"111000000000101" when"010110101010",
"111000000001000" when"010110101011",
"111000000001010" when"010110101100",
"111000000001101" when"010110101101",
"111000000010000" when"010110101110",
"111000000010011" when"010110101111",
"111000000010101" when"010110110000",
"111000000011000" when"010110110001",
"111000000011011" when"010110110010",
"111000000011101" when"010110110011",
"111000000100000" when"010110110100",
"111000000100011" when"010110110101",
"111000000100101" when"010110110110",
"111000000101000" when"010110110111",
"111000000101011" when"010110111000",
"111000000101110" when"010110111001",
"111000000110000" when"010110111010",
"111000000110011" when"010110111011",
"111000000110110" when"010110111100",
"111000000111000" when"010110111101",
"111000000111011" when"010110111110",
"111000000111110" when"010110111111",
"111000001000000" when"010111000000",
"111000001000011" when"010111000001",
"111000001000110" when"010111000010",
"111000001001000" when"010111000011",
"111000001001011" when"010111000100",
"111000001001110" when"010111000101",
"111000001010000" when"010111000110",
"111000001010011" when"010111000111",
"111000001010110" when"010111001000",
"111000001011000" when"010111001001",
"111000001011011" when"010111001010",
"111000001011110" when"010111001011",
"111000001100000" when"010111001100",
"111000001100011" when"010111001101",
"111000001100110" when"010111001110",
"111000001101000" when"010111001111",
"111000001101011" when"010111010000",
"111000001101110" when"010111010001",
"111000001110000" when"010111010010",
"111000001110011" when"010111010011",
"111000001110101" when"010111010100",
"111000001111000" when"010111010101",
"111000001111011" when"010111010110",
"111000001111101" when"010111010111",
"111000010000000" when"010111011000",
"111000010000011" when"010111011001",
"111000010000101" when"010111011010",
"111000010001000" when"010111011011",
"111000010001011" when"010111011100",
"111000010001101" when"010111011101",
"111000010010000" when"010111011110",
"111000010010010" when"010111011111",
"111000010010101" when"010111100000",
"111000010011000" when"010111100001",
"111000010011010" when"010111100010",
"111000010011101" when"010111100011",
"111000010011111" when"010111100100",
"111000010100010" when"010111100101",
"111000010100101" when"010111100110",
"111000010100111" when"010111100111",
"111000010101010" when"010111101000",
"111000010101101" when"010111101001",
"111000010101111" when"010111101010",
"111000010110010" when"010111101011",
"111000010110100" when"010111101100",
"111000010110111" when"010111101101",
"111000010111010" when"010111101110",
"111000010111100" when"010111101111",
"111000010111111" when"010111110000",
"111000011000001" when"010111110001",
"111000011000100" when"010111110010",
"111000011000110" when"010111110011",
"111000011001001" when"010111110100",
"111000011001100" when"010111110101",
"111000011001110" when"010111110110",
"111000011010001" when"010111110111",
"111000011010011" when"010111111000",
"111000011010110" when"010111111001",
"111000011011001" when"010111111010",
"111000011011011" when"010111111011",
"111000011011110" when"010111111100",
"111000011100000" when"010111111101",
"111000011100011" when"010111111110",
"111000011100101" when"010111111111",
"111000011101000" when"011000000000",
"111000011101011" when"011000000001",
"111000011101101" when"011000000010",
"111000011110000" when"011000000011",
"111000011110010" when"011000000100",
"111000011110101" when"011000000101",
"111000011110111" when"011000000110",
"111000011111010" when"011000000111",
"111000011111100" when"011000001000",
"111000011111111" when"011000001001",
"111000100000010" when"011000001010",
"111000100000100" when"011000001011",
"111000100000111" when"011000001100",
"111000100001001" when"011000001101",
"111000100001100" when"011000001110",
"111000100001110" when"011000001111",
"111000100010001" when"011000010000",
"111000100010011" when"011000010001",
"111000100010110" when"011000010010",
"111000100011000" when"011000010011",
"111000100011011" when"011000010100",
"111000100011101" when"011000010101",
"111000100100000" when"011000010110",
"111000100100011" when"011000010111",
"111000100100101" when"011000011000",
"111000100101000" when"011000011001",
"111000100101010" when"011000011010",
"111000100101101" when"011000011011",
"111000100101111" when"011000011100",
"111000100110010" when"011000011101",
"111000100110100" when"011000011110",
"111000100110111" when"011000011111",
"111000100111001" when"011000100000",
"111000100111100" when"011000100001",
"111000100111110" when"011000100010",
"111000101000001" when"011000100011",
"111000101000011" when"011000100100",
"111000101000110" when"011000100101",
"111000101001000" when"011000100110",
"111000101001011" when"011000100111",
"111000101001101" when"011000101000",
"111000101010000" when"011000101001",
"111000101010010" when"011000101010",
"111000101010101" when"011000101011",
"111000101010111" when"011000101100",
"111000101011010" when"011000101101",
"111000101011100" when"011000101110",
"111000101011111" when"011000101111",
"111000101100001" when"011000110000",
"111000101100100" when"011000110001",
"111000101100110" when"011000110010",
"111000101101001" when"011000110011",
"111000101101011" when"011000110100",
"111000101101110" when"011000110101",
"111000101110000" when"011000110110",
"111000101110011" when"011000110111",
"111000101110101" when"011000111000",
"111000101111000" when"011000111001",
"111000101111010" when"011000111010",
"111000101111100" when"011000111011",
"111000101111111" when"011000111100",
"111000110000001" when"011000111101",
"111000110000100" when"011000111110",
"111000110000110" when"011000111111",
"111000110001001" when"011001000000",
"111000110001011" when"011001000001",
"111000110001110" when"011001000010",
"111000110010000" when"011001000011",
"111000110010011" when"011001000100",
"111000110010101" when"011001000101",
"111000110011000" when"011001000110",
"111000110011010" when"011001000111",
"111000110011100" when"011001001000",
"111000110011111" when"011001001001",
"111000110100001" when"011001001010",
"111000110100100" when"011001001011",
"111000110100110" when"011001001100",
"111000110101001" when"011001001101",
"111000110101011" when"011001001110",
"111000110101110" when"011001001111",
"111000110110000" when"011001010000",
"111000110110010" when"011001010001",
"111000110110101" when"011001010010",
"111000110110111" when"011001010011",
"111000110111010" when"011001010100",
"111000110111100" when"011001010101",
"111000110111111" when"011001010110",
"111000111000001" when"011001010111",
"111000111000011" when"011001011000",
"111000111000110" when"011001011001",
"111000111001000" when"011001011010",
"111000111001011" when"011001011011",
"111000111001101" when"011001011100",
"111000111010000" when"011001011101",
"111000111010010" when"011001011110",
"111000111010100" when"011001011111",
"111000111010111" when"011001100000",
"111000111011001" when"011001100001",
"111000111011100" when"011001100010",
"111000111011110" when"011001100011",
"111000111100000" when"011001100100",
"111000111100011" when"011001100101",
"111000111100101" when"011001100110",
"111000111101000" when"011001100111",
"111000111101010" when"011001101000",
"111000111101100" when"011001101001",
"111000111101111" when"011001101010",
"111000111110001" when"011001101011",
"111000111110100" when"011001101100",
"111000111110110" when"011001101101",
"111000111111000" when"011001101110",
"111000111111011" when"011001101111",
"111000111111101" when"011001110000",
"111001000000000" when"011001110001",
"111001000000010" when"011001110010",
"111001000000100" when"011001110011",
"111001000000111" when"011001110100",
"111001000001001" when"011001110101",
"111001000001100" when"011001110110",
"111001000001110" when"011001110111",
"111001000010000" when"011001111000",
"111001000010011" when"011001111001",
"111001000010101" when"011001111010",
"111001000010111" when"011001111011",
"111001000011010" when"011001111100",
"111001000011100" when"011001111101",
"111001000011111" when"011001111110",
"111001000100001" when"011001111111",
"111001000100011" when"011010000000",
"111001000100110" when"011010000001",
"111001000101000" when"011010000010",
"111001000101010" when"011010000011",
"111001000101101" when"011010000100",
"111001000101111" when"011010000101",
"111001000110001" when"011010000110",
"111001000110100" when"011010000111",
"111001000110110" when"011010001000",
"111001000111001" when"011010001001",
"111001000111011" when"011010001010",
"111001000111101" when"011010001011",
"111001001000000" when"011010001100",
"111001001000010" when"011010001101",
"111001001000100" when"011010001110",
"111001001000111" when"011010001111",
"111001001001001" when"011010010000",
"111001001001011" when"011010010001",
"111001001001110" when"011010010010",
"111001001010000" when"011010010011",
"111001001010010" when"011010010100",
"111001001010101" when"011010010101",
"111001001010111" when"011010010110",
"111001001011001" when"011010010111",
"111001001011100" when"011010011000",
"111001001011110" when"011010011001",
"111001001100000" when"011010011010",
"111001001100011" when"011010011011",
"111001001100101" when"011010011100",
"111001001100111" when"011010011101",
"111001001101010" when"011010011110",
"111001001101100" when"011010011111",
"111001001101110" when"011010100000",
"111001001110001" when"011010100001",
"111001001110011" when"011010100010",
"111001001110101" when"011010100011",
"111001001111000" when"011010100100",
"111001001111010" when"011010100101",
"111001001111100" when"011010100110",
"111001001111111" when"011010100111",
"111001010000001" when"011010101000",
"111001010000011" when"011010101001",
"111001010000110" when"011010101010",
"111001010001000" when"011010101011",
"111001010001010" when"011010101100",
"111001010001100" when"011010101101",
"111001010001111" when"011010101110",
"111001010010001" when"011010101111",
"111001010010011" when"011010110000",
"111001010010110" when"011010110001",
"111001010011000" when"011010110010",
"111001010011010" when"011010110011",
"111001010011101" when"011010110100",
"111001010011111" when"011010110101",
"111001010100001" when"011010110110",
"111001010100011" when"011010110111",
"111001010100110" when"011010111000",
"111001010101000" when"011010111001",
"111001010101010" when"011010111010",
"111001010101101" when"011010111011",
"111001010101111" when"011010111100",
"111001010110001" when"011010111101",
"111001010110011" when"011010111110",
"111001010110110" when"011010111111",
"111001010111000" when"011011000000",
"111001010111010" when"011011000001",
"111001010111101" when"011011000010",
"111001010111111" when"011011000011",
"111001011000001" when"011011000100",
"111001011000011" when"011011000101",
"111001011000110" when"011011000110",
"111001011001000" when"011011000111",
"111001011001010" when"011011001000",
"111001011001100" when"011011001001",
"111001011001111" when"011011001010",
"111001011010001" when"011011001011",
"111001011010011" when"011011001100",
"111001011010110" when"011011001101",
"111001011011000" when"011011001110",
"111001011011010" when"011011001111",
"111001011011100" when"011011010000",
"111001011011111" when"011011010001",
"111001011100001" when"011011010010",
"111001011100011" when"011011010011",
"111001011100101" when"011011010100",
"111001011101000" when"011011010101",
"111001011101010" when"011011010110",
"111001011101100" when"011011010111",
"111001011101110" when"011011011000",
"111001011110001" when"011011011001",
"111001011110011" when"011011011010",
"111001011110101" when"011011011011",
"111001011110111" when"011011011100",
"111001011111010" when"011011011101",
"111001011111100" when"011011011110",
"111001011111110" when"011011011111",
"111001100000000" when"011011100000",
"111001100000011" when"011011100001",
"111001100000101" when"011011100010",
"111001100000111" when"011011100011",
"111001100001001" when"011011100100",
"111001100001011" when"011011100101",
"111001100001110" when"011011100110",
"111001100010000" when"011011100111",
"111001100010010" when"011011101000",
"111001100010100" when"011011101001",
"111001100010111" when"011011101010",
"111001100011001" when"011011101011",
"111001100011011" when"011011101100",
"111001100011101" when"011011101101",
"111001100011111" when"011011101110",
"111001100100010" when"011011101111",
"111001100100100" when"011011110000",
"111001100100110" when"011011110001",
"111001100101000" when"011011110010",
"111001100101011" when"011011110011",
"111001100101101" when"011011110100",
"111001100101111" when"011011110101",
"111001100110001" when"011011110110",
"111001100110011" when"011011110111",
"111001100110110" when"011011111000",
"111001100111000" when"011011111001",
"111001100111010" when"011011111010",
"111001100111100" when"011011111011",
"111001100111110" when"011011111100",
"111001101000001" when"011011111101",
"111001101000011" when"011011111110",
"111001101000101" when"011011111111",
"111001101000111" when"011100000000",
"111001101001001" when"011100000001",
"111001101001100" when"011100000010",
"111001101001110" when"011100000011",
"111001101010000" when"011100000100",
"111001101010010" when"011100000101",
"111001101010100" when"011100000110",
"111001101010111" when"011100000111",
"111001101011001" when"011100001000",
"111001101011011" when"011100001001",
"111001101011101" when"011100001010",
"111001101011111" when"011100001011",
"111001101100010" when"011100001100",
"111001101100100" when"011100001101",
"111001101100110" when"011100001110",
"111001101101000" when"011100001111",
"111001101101010" when"011100010000",
"111001101101100" when"011100010001",
"111001101101111" when"011100010010",
"111001101110001" when"011100010011",
"111001101110011" when"011100010100",
"111001101110101" when"011100010101",
"111001101110111" when"011100010110",
"111001101111001" when"011100010111",
"111001101111100" when"011100011000",
"111001101111110" when"011100011001",
"111001110000000" when"011100011010",
"111001110000010" when"011100011011",
"111001110000100" when"011100011100",
"111001110000110" when"011100011101",
"111001110001001" when"011100011110",
"111001110001011" when"011100011111",
"111001110001101" when"011100100000",
"111001110001111" when"011100100001",
"111001110010001" when"011100100010",
"111001110010011" when"011100100011",
"111001110010110" when"011100100100",
"111001110011000" when"011100100101",
"111001110011010" when"011100100110",
"111001110011100" when"011100100111",
"111001110011110" when"011100101000",
"111001110100000" when"011100101001",
"111001110100011" when"011100101010",
"111001110100101" when"011100101011",
"111001110100111" when"011100101100",
"111001110101001" when"011100101101",
"111001110101011" when"011100101110",
"111001110101101" when"011100101111",
"111001110101111" when"011100110000",
"111001110110010" when"011100110001",
"111001110110100" when"011100110010",
"111001110110110" when"011100110011",
"111001110111000" when"011100110100",
"111001110111010" when"011100110101",
"111001110111100" when"011100110110",
"111001110111110" when"011100110111",
"111001111000000" when"011100111000",
"111001111000011" when"011100111001",
"111001111000101" when"011100111010",
"111001111000111" when"011100111011",
"111001111001001" when"011100111100",
"111001111001011" when"011100111101",
"111001111001101" when"011100111110",
"111001111001111" when"011100111111",
"111001111010001" when"011101000000",
"111001111010100" when"011101000001",
"111001111010110" when"011101000010",
"111001111011000" when"011101000011",
"111001111011010" when"011101000100",
"111001111011100" when"011101000101",
"111001111011110" when"011101000110",
"111001111100000" when"011101000111",
"111001111100010" when"011101001000",
"111001111100101" when"011101001001",
"111001111100111" when"011101001010",
"111001111101001" when"011101001011",
"111001111101011" when"011101001100",
"111001111101101" when"011101001101",
"111001111101111" when"011101001110",
"111001111110001" when"011101001111",
"111001111110011" when"011101010000",
"111001111110101" when"011101010001",
"111001111111000" when"011101010010",
"111001111111010" when"011101010011",
"111001111111100" when"011101010100",
"111001111111110" when"011101010101",
"111010000000000" when"011101010110",
"111010000000010" when"011101010111",
"111010000000100" when"011101011000",
"111010000000110" when"011101011001",
"111010000001000" when"011101011010",
"111010000001010" when"011101011011",
"111010000001100" when"011101011100",
"111010000001111" when"011101011101",
"111010000010001" when"011101011110",
"111010000010011" when"011101011111",
"111010000010101" when"011101100000",
"111010000010111" when"011101100001",
"111010000011001" when"011101100010",
"111010000011011" when"011101100011",
"111010000011101" when"011101100100",
"111010000011111" when"011101100101",
"111010000100001" when"011101100110",
"111010000100011" when"011101100111",
"111010000100101" when"011101101000",
"111010000101000" when"011101101001",
"111010000101010" when"011101101010",
"111010000101100" when"011101101011",
"111010000101110" when"011101101100",
"111010000110000" when"011101101101",
"111010000110010" when"011101101110",
"111010000110100" when"011101101111",
"111010000110110" when"011101110000",
"111010000111000" when"011101110001",
"111010000111010" when"011101110010",
"111010000111100" when"011101110011",
"111010000111110" when"011101110100",
"111010001000000" when"011101110101",
"111010001000010" when"011101110110",
"111010001000101" when"011101110111",
"111010001000111" when"011101111000",
"111010001001001" when"011101111001",
"111010001001011" when"011101111010",
"111010001001101" when"011101111011",
"111010001001111" when"011101111100",
"111010001010001" when"011101111101",
"111010001010011" when"011101111110",
"111010001010101" when"011101111111",
"111010001010111" when"011110000000",
"111010001011001" when"011110000001",
"111010001011011" when"011110000010",
"111010001011101" when"011110000011",
"111010001011111" when"011110000100",
"111010001100001" when"011110000101",
"111010001100011" when"011110000110",
"111010001100101" when"011110000111",
"111010001100111" when"011110001000",
"111010001101001" when"011110001001",
"111010001101100" when"011110001010",
"111010001101110" when"011110001011",
"111010001110000" when"011110001100",
"111010001110010" when"011110001101",
"111010001110100" when"011110001110",
"111010001110110" when"011110001111",
"111010001111000" when"011110010000",
"111010001111010" when"011110010001",
"111010001111100" when"011110010010",
"111010001111110" when"011110010011",
"111010010000000" when"011110010100",
"111010010000010" when"011110010101",
"111010010000100" when"011110010110",
"111010010000110" when"011110010111",
"111010010001000" when"011110011000",
"111010010001010" when"011110011001",
"111010010001100" when"011110011010",
"111010010001110" when"011110011011",
"111010010010000" when"011110011100",
"111010010010010" when"011110011101",
"111010010010100" when"011110011110",
"111010010010110" when"011110011111",
"111010010011000" when"011110100000",
"111010010011010" when"011110100001",
"111010010011100" when"011110100010",
"111010010011110" when"011110100011",
"111010010100000" when"011110100100",
"111010010100010" when"011110100101",
"111010010100100" when"011110100110",
"111010010100110" when"011110100111",
"111010010101000" when"011110101000",
"111010010101010" when"011110101001",
"111010010101100" when"011110101010",
"111010010101110" when"011110101011",
"111010010110000" when"011110101100",
"111010010110010" when"011110101101",
"111010010110100" when"011110101110",
"111010010110110" when"011110101111",
"111010010111000" when"011110110000",
"111010010111010" when"011110110001",
"111010010111100" when"011110110010",
"111010010111110" when"011110110011",
"111010011000000" when"011110110100",
"111010011000010" when"011110110101",
"111010011000100" when"011110110110",
"111010011000110" when"011110110111",
"111010011001000" when"011110111000",
"111010011001010" when"011110111001",
"111010011001100" when"011110111010",
"111010011001110" when"011110111011",
"111010011010000" when"011110111100",
"111010011010010" when"011110111101",
"111010011010100" when"011110111110",
"111010011010110" when"011110111111",
"111010011011000" when"011111000000",
"111010011011010" when"011111000001",
"111010011011100" when"011111000010",
"111010011011110" when"011111000011",
"111010011100000" when"011111000100",
"111010011100010" when"011111000101",
"111010011100100" when"011111000110",
"111010011100110" when"011111000111",
"111010011101000" when"011111001000",
"111010011101010" when"011111001001",
"111010011101100" when"011111001010",
"111010011101110" when"011111001011",
"111010011110000" when"011111001100",
"111010011110010" when"011111001101",
"111010011110100" when"011111001110",
"111010011110110" when"011111001111",
"111010011111000" when"011111010000",
"111010011111010" when"011111010001",
"111010011111100" when"011111010010",
"111010011111110" when"011111010011",
"111010100000000" when"011111010100",
"111010100000010" when"011111010101",
"111010100000100" when"011111010110",
"111010100000110" when"011111010111",
"111010100001000" when"011111011000",
"111010100001010" when"011111011001",
"111010100001100" when"011111011010",
"111010100001101" when"011111011011",
"111010100001111" when"011111011100",
"111010100010001" when"011111011101",
"111010100010011" when"011111011110",
"111010100010101" when"011111011111",
"111010100010111" when"011111100000",
"111010100011001" when"011111100001",
"111010100011011" when"011111100010",
"111010100011101" when"011111100011",
"111010100011111" when"011111100100",
"111010100100001" when"011111100101",
"111010100100011" when"011111100110",
"111010100100101" when"011111100111",
"111010100100111" when"011111101000",
"111010100101001" when"011111101001",
"111010100101011" when"011111101010",
"111010100101101" when"011111101011",
"111010100101111" when"011111101100",
"111010100110001" when"011111101101",
"111010100110011" when"011111101110",
"111010100110100" when"011111101111",
"111010100110110" when"011111110000",
"111010100111000" when"011111110001",
"111010100111010" when"011111110010",
"111010100111100" when"011111110011",
"111010100111110" when"011111110100",
"111010101000000" when"011111110101",
"111010101000010" when"011111110110",
"111010101000100" when"011111110111",
"111010101000110" when"011111111000",
"111010101001000" when"011111111001",
"111010101001010" when"011111111010",
"111010101001100" when"011111111011",
"111010101001110" when"011111111100",
"111010101010000" when"011111111101",
"111010101010001" when"011111111110",
"111010101010011" when"011111111111",
"111010101010101" when"100000000000",
"111010101010111" when"100000000001",
"111010101011001" when"100000000010",
"111010101011011" when"100000000011",
"111010101011101" when"100000000100",
"111010101011111" when"100000000101",
"111010101100001" when"100000000110",
"111010101100011" when"100000000111",
"111010101100101" when"100000001000",
"111010101100111" when"100000001001",
"111010101101000" when"100000001010",
"111010101101010" when"100000001011",
"111010101101100" when"100000001100",
"111010101101110" when"100000001101",
"111010101110000" when"100000001110",
"111010101110010" when"100000001111",
"111010101110100" when"100000010000",
"111010101110110" when"100000010001",
"111010101111000" when"100000010010",
"111010101111010" when"100000010011",
"111010101111100" when"100000010100",
"111010101111101" when"100000010101",
"111010101111111" when"100000010110",
"111010110000001" when"100000010111",
"111010110000011" when"100000011000",
"111010110000101" when"100000011001",
"111010110000111" when"100000011010",
"111010110001001" when"100000011011",
"111010110001011" when"100000011100",
"111010110001101" when"100000011101",
"111010110001111" when"100000011110",
"111010110010000" when"100000011111",
"111010110010010" when"100000100000",
"111010110010100" when"100000100001",
"111010110010110" when"100000100010",
"111010110011000" when"100000100011",
"111010110011010" when"100000100100",
"111010110011100" when"100000100101",
"111010110011110" when"100000100110",
"111010110100000" when"100000100111",
"111010110100010" when"100000101000",
"111010110100011" when"100000101001",
"111010110100101" when"100000101010",
"111010110100111" when"100000101011",
"111010110101001" when"100000101100",
"111010110101011" when"100000101101",
"111010110101101" when"100000101110",
"111010110101111" when"100000101111",
"111010110110001" when"100000110000",
"111010110110010" when"100000110001",
"111010110110100" when"100000110010",
"111010110110110" when"100000110011",
"111010110111000" when"100000110100",
"111010110111010" when"100000110101",
"111010110111100" when"100000110110",
"111010110111110" when"100000110111",
"111010111000000" when"100000111000",
"111010111000001" when"100000111001",
"111010111000011" when"100000111010",
"111010111000101" when"100000111011",
"111010111000111" when"100000111100",
"111010111001001" when"100000111101",
"111010111001011" when"100000111110",
"111010111001101" when"100000111111",
"111010111001111" when"100001000000",
"111010111010000" when"100001000001",
"111010111010010" when"100001000010",
"111010111010100" when"100001000011",
"111010111010110" when"100001000100",
"111010111011000" when"100001000101",
"111010111011010" when"100001000110",
"111010111011100" when"100001000111",
"111010111011101" when"100001001000",
"111010111011111" when"100001001001",
"111010111100001" when"100001001010",
"111010111100011" when"100001001011",
"111010111100101" when"100001001100",
"111010111100111" when"100001001101",
"111010111101001" when"100001001110",
"111010111101010" when"100001001111",
"111010111101100" when"100001010000",
"111010111101110" when"100001010001",
"111010111110000" when"100001010010",
"111010111110010" when"100001010011",
"111010111110100" when"100001010100",
"111010111110110" when"100001010101",
"111010111110111" when"100001010110",
"111010111111001" when"100001010111",
"111010111111011" when"100001011000",
"111010111111101" when"100001011001",
"111010111111111" when"100001011010",
"111011000000001" when"100001011011",
"111011000000010" when"100001011100",
"111011000000100" when"100001011101",
"111011000000110" when"100001011110",
"111011000001000" when"100001011111",
"111011000001010" when"100001100000",
"111011000001100" when"100001100001",
"111011000001101" when"100001100010",
"111011000001111" when"100001100011",
"111011000010001" when"100001100100",
"111011000010011" when"100001100101",
"111011000010101" when"100001100110",
"111011000010111" when"100001100111",
"111011000011000" when"100001101000",
"111011000011010" when"100001101001",
"111011000011100" when"100001101010",
"111011000011110" when"100001101011",
"111011000100000" when"100001101100",
"111011000100010" when"100001101101",
"111011000100011" when"100001101110",
"111011000100101" when"100001101111",
"111011000100111" when"100001110000",
"111011000101001" when"100001110001",
"111011000101011" when"100001110010",
"111011000101101" when"100001110011",
"111011000101110" when"100001110100",
"111011000110000" when"100001110101",
"111011000110010" when"100001110110",
"111011000110100" when"100001110111",
"111011000110110" when"100001111000",
"111011000110111" when"100001111001",
"111011000111001" when"100001111010",
"111011000111011" when"100001111011",
"111011000111101" when"100001111100",
"111011000111111" when"100001111101",
"111011001000001" when"100001111110",
"111011001000010" when"100001111111",
"111011001000100" when"100010000000",
"111011001000110" when"100010000001",
"111011001001000" when"100010000010",
"111011001001010" when"100010000011",
"111011001001011" when"100010000100",
"111011001001101" when"100010000101",
"111011001001111" when"100010000110",
"111011001010001" when"100010000111",
"111011001010011" when"100010001000",
"111011001010100" when"100010001001",
"111011001010110" when"100010001010",
"111011001011000" when"100010001011",
"111011001011010" when"100010001100",
"111011001011100" when"100010001101",
"111011001011101" when"100010001110",
"111011001011111" when"100010001111",
"111011001100001" when"100010010000",
"111011001100011" when"100010010001",
"111011001100101" when"100010010010",
"111011001100110" when"100010010011",
"111011001101000" when"100010010100",
"111011001101010" when"100010010101",
"111011001101100" when"100010010110",
"111011001101110" when"100010010111",
"111011001101111" when"100010011000",
"111011001110001" when"100010011001",
"111011001110011" when"100010011010",
"111011001110101" when"100010011011",
"111011001110110" when"100010011100",
"111011001111000" when"100010011101",
"111011001111010" when"100010011110",
"111011001111100" when"100010011111",
"111011001111110" when"100010100000",
"111011001111111" when"100010100001",
"111011010000001" when"100010100010",
"111011010000011" when"100010100011",
"111011010000101" when"100010100100",
"111011010000111" when"100010100101",
"111011010001000" when"100010100110",
"111011010001010" when"100010100111",
"111011010001100" when"100010101000",
"111011010001110" when"100010101001",
"111011010001111" when"100010101010",
"111011010010001" when"100010101011",
"111011010010011" when"100010101100",
"111011010010101" when"100010101101",
"111011010010111" when"100010101110",
"111011010011000" when"100010101111",
"111011010011010" when"100010110000",
"111011010011100" when"100010110001",
"111011010011110" when"100010110010",
"111011010011111" when"100010110011",
"111011010100001" when"100010110100",
"111011010100011" when"100010110101",
"111011010100101" when"100010110110",
"111011010100110" when"100010110111",
"111011010101000" when"100010111000",
"111011010101010" when"100010111001",
"111011010101100" when"100010111010",
"111011010101110" when"100010111011",
"111011010101111" when"100010111100",
"111011010110001" when"100010111101",
"111011010110011" when"100010111110",
"111011010110101" when"100010111111",
"111011010110110" when"100011000000",
"111011010111000" when"100011000001",
"111011010111010" when"100011000010",
"111011010111100" when"100011000011",
"111011010111101" when"100011000100",
"111011010111111" when"100011000101",
"111011011000001" when"100011000110",
"111011011000011" when"100011000111",
"111011011000100" when"100011001000",
"111011011000110" when"100011001001",
"111011011001000" when"100011001010",
"111011011001010" when"100011001011",
"111011011001011" when"100011001100",
"111011011001101" when"100011001101",
"111011011001111" when"100011001110",
"111011011010001" when"100011001111",
"111011011010010" when"100011010000",
"111011011010100" when"100011010001",
"111011011010110" when"100011010010",
"111011011011000" when"100011010011",
"111011011011001" when"100011010100",
"111011011011011" when"100011010101",
"111011011011101" when"100011010110",
"111011011011111" when"100011010111",
"111011011100000" when"100011011000",
"111011011100010" when"100011011001",
"111011011100100" when"100011011010",
"111011011100110" when"100011011011",
"111011011100111" when"100011011100",
"111011011101001" when"100011011101",
"111011011101011" when"100011011110",
"111011011101100" when"100011011111",
"111011011101110" when"100011100000",
"111011011110000" when"100011100001",
"111011011110010" when"100011100010",
"111011011110011" when"100011100011",
"111011011110101" when"100011100100",
"111011011110111" when"100011100101",
"111011011111001" when"100011100110",
"111011011111010" when"100011100111",
"111011011111100" when"100011101000",
"111011011111110" when"100011101001",
"111011100000000" when"100011101010",
"111011100000001" when"100011101011",
"111011100000011" when"100011101100",
"111011100000101" when"100011101101",
"111011100000110" when"100011101110",
"111011100001000" when"100011101111",
"111011100001010" when"100011110000",
"111011100001100" when"100011110001",
"111011100001101" when"100011110010",
"111011100001111" when"100011110011",
"111011100010001" when"100011110100",
"111011100010010" when"100011110101",
"111011100010100" when"100011110110",
"111011100010110" when"100011110111",
"111011100011000" when"100011111000",
"111011100011001" when"100011111001",
"111011100011011" when"100011111010",
"111011100011101" when"100011111011",
"111011100011110" when"100011111100",
"111011100100000" when"100011111101",
"111011100100010" when"100011111110",
"111011100100100" when"100011111111",
"111011100100101" when"100100000000",
"111011100100111" when"100100000001",
"111011100101001" when"100100000010",
"111011100101010" when"100100000011",
"111011100101100" when"100100000100",
"111011100101110" when"100100000101",
"111011100110000" when"100100000110",
"111011100110001" when"100100000111",
"111011100110011" when"100100001000",
"111011100110101" when"100100001001",
"111011100110110" when"100100001010",
"111011100111000" when"100100001011",
"111011100111010" when"100100001100",
"111011100111011" when"100100001101",
"111011100111101" when"100100001110",
"111011100111111" when"100100001111",
"111011101000001" when"100100010000",
"111011101000010" when"100100010001",
"111011101000100" when"100100010010",
"111011101000110" when"100100010011",
"111011101000111" when"100100010100",
"111011101001001" when"100100010101",
"111011101001011" when"100100010110",
"111011101001100" when"100100010111",
"111011101001110" when"100100011000",
"111011101010000" when"100100011001",
"111011101010010" when"100100011010",
"111011101010011" when"100100011011",
"111011101010101" when"100100011100",
"111011101010111" when"100100011101",
"111011101011000" when"100100011110",
"111011101011010" when"100100011111",
"111011101011100" when"100100100000",
"111011101011101" when"100100100001",
"111011101011111" when"100100100010",
"111011101100001" when"100100100011",
"111011101100010" when"100100100100",
"111011101100100" when"100100100101",
"111011101100110" when"100100100110",
"111011101100111" when"100100100111",
"111011101101001" when"100100101000",
"111011101101011" when"100100101001",
"111011101101100" when"100100101010",
"111011101101110" when"100100101011",
"111011101110000" when"100100101100",
"111011101110010" when"100100101101",
"111011101110011" when"100100101110",
"111011101110101" when"100100101111",
"111011101110111" when"100100110000",
"111011101111000" when"100100110001",
"111011101111010" when"100100110010",
"111011101111100" when"100100110011",
"111011101111101" when"100100110100",
"111011101111111" when"100100110101",
"111011110000001" when"100100110110",
"111011110000010" when"100100110111",
"111011110000100" when"100100111000",
"111011110000110" when"100100111001",
"111011110000111" when"100100111010",
"111011110001001" when"100100111011",
"111011110001011" when"100100111100",
"111011110001100" when"100100111101",
"111011110001110" when"100100111110",
"111011110010000" when"100100111111",
"111011110010001" when"100101000000",
"111011110010011" when"100101000001",
"111011110010101" when"100101000010",
"111011110010110" when"100101000011",
"111011110011000" when"100101000100",
"111011110011010" when"100101000101",
"111011110011011" when"100101000110",
"111011110011101" when"100101000111",
"111011110011111" when"100101001000",
"111011110100000" when"100101001001",
"111011110100010" when"100101001010",
"111011110100100" when"100101001011",
"111011110100101" when"100101001100",
"111011110100111" when"100101001101",
"111011110101000" when"100101001110",
"111011110101010" when"100101001111",
"111011110101100" when"100101010000",
"111011110101101" when"100101010001",
"111011110101111" when"100101010010",
"111011110110001" when"100101010011",
"111011110110010" when"100101010100",
"111011110110100" when"100101010101",
"111011110110110" when"100101010110",
"111011110110111" when"100101010111",
"111011110111001" when"100101011000",
"111011110111011" when"100101011001",
"111011110111100" when"100101011010",
"111011110111110" when"100101011011",
"111011111000000" when"100101011100",
"111011111000001" when"100101011101",
"111011111000011" when"100101011110",
"111011111000100" when"100101011111",
"111011111000110" when"100101100000",
"111011111001000" when"100101100001",
"111011111001001" when"100101100010",
"111011111001011" when"100101100011",
"111011111001101" when"100101100100",
"111011111001110" when"100101100101",
"111011111010000" when"100101100110",
"111011111010010" when"100101100111",
"111011111010011" when"100101101000",
"111011111010101" when"100101101001",
"111011111010111" when"100101101010",
"111011111011000" when"100101101011",
"111011111011010" when"100101101100",
"111011111011011" when"100101101101",
"111011111011101" when"100101101110",
"111011111011111" when"100101101111",
"111011111100000" when"100101110000",
"111011111100010" when"100101110001",
"111011111100100" when"100101110010",
"111011111100101" when"100101110011",
"111011111100111" when"100101110100",
"111011111101000" when"100101110101",
"111011111101010" when"100101110110",
"111011111101100" when"100101110111",
"111011111101101" when"100101111000",
"111011111101111" when"100101111001",
"111011111110001" when"100101111010",
"111011111110010" when"100101111011",
"111011111110100" when"100101111100",
"111011111110101" when"100101111101",
"111011111110111" when"100101111110",
"111011111111001" when"100101111111",
"111011111111010" when"100110000000",
"111011111111100" when"100110000001",
"111011111111110" when"100110000010",
"111011111111111" when"100110000011",
"111100000000001" when"100110000100",
"111100000000010" when"100110000101",
"111100000000100" when"100110000110",
"111100000000110" when"100110000111",
"111100000000111" when"100110001000",
"111100000001001" when"100110001001",
"111100000001010" when"100110001010",
"111100000001100" when"100110001011",
"111100000001110" when"100110001100",
"111100000001111" when"100110001101",
"111100000010001" when"100110001110",
"111100000010011" when"100110001111",
"111100000010100" when"100110010000",
"111100000010110" when"100110010001",
"111100000010111" when"100110010010",
"111100000011001" when"100110010011",
"111100000011011" when"100110010100",
"111100000011100" when"100110010101",
"111100000011110" when"100110010110",
"111100000011111" when"100110010111",
"111100000100001" when"100110011000",
"111100000100011" when"100110011001",
"111100000100100" when"100110011010",
"111100000100110" when"100110011011",
"111100000100111" when"100110011100",
"111100000101001" when"100110011101",
"111100000101011" when"100110011110",
"111100000101100" when"100110011111",
"111100000101110" when"100110100000",
"111100000101111" when"100110100001",
"111100000110001" when"100110100010",
"111100000110011" when"100110100011",
"111100000110100" when"100110100100",
"111100000110110" when"100110100101",
"111100000110111" when"100110100110",
"111100000111001" when"100110100111",
"111100000111011" when"100110101000",
"111100000111100" when"100110101001",
"111100000111110" when"100110101010",
"111100000111111" when"100110101011",
"111100001000001" when"100110101100",
"111100001000011" when"100110101101",
"111100001000100" when"100110101110",
"111100001000110" when"100110101111",
"111100001000111" when"100110110000",
"111100001001001" when"100110110001",
"111100001001010" when"100110110010",
"111100001001100" when"100110110011",
"111100001001110" when"100110110100",
"111100001001111" when"100110110101",
"111100001010001" when"100110110110",
"111100001010010" when"100110110111",
"111100001010100" when"100110111000",
"111100001010110" when"100110111001",
"111100001010111" when"100110111010",
"111100001011001" when"100110111011",
"111100001011010" when"100110111100",
"111100001011100" when"100110111101",
"111100001011101" when"100110111110",
"111100001011111" when"100110111111",
"111100001100001" when"100111000000",
"111100001100010" when"100111000001",
"111100001100100" when"100111000010",
"111100001100101" when"100111000011",
"111100001100111" when"100111000100",
"111100001101001" when"100111000101",
"111100001101010" when"100111000110",
"111100001101100" when"100111000111",
"111100001101101" when"100111001000",
"111100001101111" when"100111001001",
"111100001110000" when"100111001010",
"111100001110010" when"100111001011",
"111100001110100" when"100111001100",
"111100001110101" when"100111001101",
"111100001110111" when"100111001110",
"111100001111000" when"100111001111",
"111100001111010" when"100111010000",
"111100001111011" when"100111010001",
"111100001111101" when"100111010010",
"111100001111111" when"100111010011",
"111100010000000" when"100111010100",
"111100010000010" when"100111010101",
"111100010000011" when"100111010110",
"111100010000101" when"100111010111",
"111100010000110" when"100111011000",
"111100010001000" when"100111011001",
"111100010001001" when"100111011010",
"111100010001011" when"100111011011",
"111100010001101" when"100111011100",
"111100010001110" when"100111011101",
"111100010010000" when"100111011110",
"111100010010001" when"100111011111",
"111100010010011" when"100111100000",
"111100010010100" when"100111100001",
"111100010010110" when"100111100010",
"111100010010111" when"100111100011",
"111100010011001" when"100111100100",
"111100010011011" when"100111100101",
"111100010011100" when"100111100110",
"111100010011110" when"100111100111",
"111100010011111" when"100111101000",
"111100010100001" when"100111101001",
"111100010100010" when"100111101010",
"111100010100100" when"100111101011",
"111100010100101" when"100111101100",
"111100010100111" when"100111101101",
"111100010101001" when"100111101110",
"111100010101010" when"100111101111",
"111100010101100" when"100111110000",
"111100010101101" when"100111110001",
"111100010101111" when"100111110010",
"111100010110000" when"100111110011",
"111100010110010" when"100111110100",
"111100010110011" when"100111110101",
"111100010110101" when"100111110110",
"111100010110111" when"100111110111",
"111100010111000" when"100111111000",
"111100010111010" when"100111111001",
"111100010111011" when"100111111010",
"111100010111101" when"100111111011",
"111100010111110" when"100111111100",
"111100011000000" when"100111111101",
"111100011000001" when"100111111110",
"111100011000011" when"100111111111",
"111100011000100" when"101000000000",
"111100011000110" when"101000000001",
"111100011000111" when"101000000010",
"111100011001001" when"101000000011",
"111100011001011" when"101000000100",
"111100011001100" when"101000000101",
"111100011001110" when"101000000110",
"111100011001111" when"101000000111",
"111100011010001" when"101000001000",
"111100011010010" when"101000001001",
"111100011010100" when"101000001010",
"111100011010101" when"101000001011",
"111100011010111" when"101000001100",
"111100011011000" when"101000001101",
"111100011011010" when"101000001110",
"111100011011011" when"101000001111",
"111100011011101" when"101000010000",
"111100011011110" when"101000010001",
"111100011100000" when"101000010010",
"111100011100010" when"101000010011",
"111100011100011" when"101000010100",
"111100011100101" when"101000010101",
"111100011100110" when"101000010110",
"111100011101000" when"101000010111",
"111100011101001" when"101000011000",
"111100011101011" when"101000011001",
"111100011101100" when"101000011010",
"111100011101110" when"101000011011",
"111100011101111" when"101000011100",
"111100011110001" when"101000011101",
"111100011110010" when"101000011110",
"111100011110100" when"101000011111",
"111100011110101" when"101000100000",
"111100011110111" when"101000100001",
"111100011111000" when"101000100010",
"111100011111010" when"101000100011",
"111100011111011" when"101000100100",
"111100011111101" when"101000100101",
"111100011111110" when"101000100110",
"111100100000000" when"101000100111",
"111100100000001" when"101000101000",
"111100100000011" when"101000101001",
"111100100000100" when"101000101010",
"111100100000110" when"101000101011",
"111100100001000" when"101000101100",
"111100100001001" when"101000101101",
"111100100001011" when"101000101110",
"111100100001100" when"101000101111",
"111100100001110" when"101000110000",
"111100100001111" when"101000110001",
"111100100010001" when"101000110010",
"111100100010010" when"101000110011",
"111100100010100" when"101000110100",
"111100100010101" when"101000110101",
"111100100010111" when"101000110110",
"111100100011000" when"101000110111",
"111100100011010" when"101000111000",
"111100100011011" when"101000111001",
"111100100011101" when"101000111010",
"111100100011110" when"101000111011",
"111100100100000" when"101000111100",
"111100100100001" when"101000111101",
"111100100100011" when"101000111110",
"111100100100100" when"101000111111",
"111100100100110" when"101001000000",
"111100100100111" when"101001000001",
"111100100101001" when"101001000010",
"111100100101010" when"101001000011",
"111100100101100" when"101001000100",
"111100100101101" when"101001000101",
"111100100101111" when"101001000110",
"111100100110000" when"101001000111",
"111100100110010" when"101001001000",
"111100100110011" when"101001001001",
"111100100110101" when"101001001010",
"111100100110110" when"101001001011",
"111100100111000" when"101001001100",
"111100100111001" when"101001001101",
"111100100111011" when"101001001110",
"111100100111100" when"101001001111",
"111100100111110" when"101001010000",
"111100100111111" when"101001010001",
"111100101000001" when"101001010010",
"111100101000010" when"101001010011",
"111100101000100" when"101001010100",
"111100101000101" when"101001010101",
"111100101000111" when"101001010110",
"111100101001000" when"101001010111",
"111100101001010" when"101001011000",
"111100101001011" when"101001011001",
"111100101001100" when"101001011010",
"111100101001110" when"101001011011",
"111100101001111" when"101001011100",
"111100101010001" when"101001011101",
"111100101010010" when"101001011110",
"111100101010100" when"101001011111",
"111100101010101" when"101001100000",
"111100101010111" when"101001100001",
"111100101011000" when"101001100010",
"111100101011010" when"101001100011",
"111100101011011" when"101001100100",
"111100101011101" when"101001100101",
"111100101011110" when"101001100110",
"111100101100000" when"101001100111",
"111100101100001" when"101001101000",
"111100101100011" when"101001101001",
"111100101100100" when"101001101010",
"111100101100110" when"101001101011",
"111100101100111" when"101001101100",
"111100101101001" when"101001101101",
"111100101101010" when"101001101110",
"111100101101100" when"101001101111",
"111100101101101" when"101001110000",
"111100101101111" when"101001110001",
"111100101110000" when"101001110010",
"111100101110001" when"101001110011",
"111100101110011" when"101001110100",
"111100101110100" when"101001110101",
"111100101110110" when"101001110110",
"111100101110111" when"101001110111",
"111100101111001" when"101001111000",
"111100101111010" when"101001111001",
"111100101111100" when"101001111010",
"111100101111101" when"101001111011",
"111100101111111" when"101001111100",
"111100110000000" when"101001111101",
"111100110000010" when"101001111110",
"111100110000011" when"101001111111",
"111100110000101" when"101010000000",
"111100110000110" when"101010000001",
"111100110001000" when"101010000010",
"111100110001001" when"101010000011",
"111100110001010" when"101010000100",
"111100110001100" when"101010000101",
"111100110001101" when"101010000110",
"111100110001111" when"101010000111",
"111100110010000" when"101010001000",
"111100110010010" when"101010001001",
"111100110010011" when"101010001010",
"111100110010101" when"101010001011",
"111100110010110" when"101010001100",
"111100110011000" when"101010001101",
"111100110011001" when"101010001110",
"111100110011011" when"101010001111",
"111100110011100" when"101010010000",
"111100110011101" when"101010010001",
"111100110011111" when"101010010010",
"111100110100000" when"101010010011",
"111100110100010" when"101010010100",
"111100110100011" when"101010010101",
"111100110100101" when"101010010110",
"111100110100110" when"101010010111",
"111100110101000" when"101010011000",
"111100110101001" when"101010011001",
"111100110101011" when"101010011010",
"111100110101100" when"101010011011",
"111100110101101" when"101010011100",
"111100110101111" when"101010011101",
"111100110110000" when"101010011110",
"111100110110010" when"101010011111",
"111100110110011" when"101010100000",
"111100110110101" when"101010100001",
"111100110110110" when"101010100010",
"111100110111000" when"101010100011",
"111100110111001" when"101010100100",
"111100110111010" when"101010100101",
"111100110111100" when"101010100110",
"111100110111101" when"101010100111",
"111100110111111" when"101010101000",
"111100111000000" when"101010101001",
"111100111000010" when"101010101010",
"111100111000011" when"101010101011",
"111100111000101" when"101010101100",
"111100111000110" when"101010101101",
"111100111000111" when"101010101110",
"111100111001001" when"101010101111",
"111100111001010" when"101010110000",
"111100111001100" when"101010110001",
"111100111001101" when"101010110010",
"111100111001111" when"101010110011",
"111100111010000" when"101010110100",
"111100111010010" when"101010110101",
"111100111010011" when"101010110110",
"111100111010100" when"101010110111",
"111100111010110" when"101010111000",
"111100111010111" when"101010111001",
"111100111011001" when"101010111010",
"111100111011010" when"101010111011",
"111100111011100" when"101010111100",
"111100111011101" when"101010111101",
"111100111011110" when"101010111110",
"111100111100000" when"101010111111",
"111100111100001" when"101011000000",
"111100111100011" when"101011000001",
"111100111100100" when"101011000010",
"111100111100110" when"101011000011",
"111100111100111" when"101011000100",
"111100111101000" when"101011000101",
"111100111101010" when"101011000110",
"111100111101011" when"101011000111",
"111100111101101" when"101011001000",
"111100111101110" when"101011001001",
"111100111110000" when"101011001010",
"111100111110001" when"101011001011",
"111100111110010" when"101011001100",
"111100111110100" when"101011001101",
"111100111110101" when"101011001110",
"111100111110111" when"101011001111",
"111100111111000" when"101011010000",
"111100111111010" when"101011010001",
"111100111111011" when"101011010010",
"111100111111100" when"101011010011",
"111100111111110" when"101011010100",
"111100111111111" when"101011010101",
"111101000000001" when"101011010110",
"111101000000010" when"101011010111",
"111101000000011" when"101011011000",
"111101000000101" when"101011011001",
"111101000000110" when"101011011010",
"111101000001000" when"101011011011",
"111101000001001" when"101011011100",
"111101000001011" when"101011011101",
"111101000001100" when"101011011110",
"111101000001101" when"101011011111",
"111101000001111" when"101011100000",
"111101000010000" when"101011100001",
"111101000010010" when"101011100010",
"111101000010011" when"101011100011",
"111101000010100" when"101011100100",
"111101000010110" when"101011100101",
"111101000010111" when"101011100110",
"111101000011001" when"101011100111",
"111101000011010" when"101011101000",
"111101000011100" when"101011101001",
"111101000011101" when"101011101010",
"111101000011110" when"101011101011",
"111101000100000" when"101011101100",
"111101000100001" when"101011101101",
"111101000100011" when"101011101110",
"111101000100100" when"101011101111",
"111101000100101" when"101011110000",
"111101000100111" when"101011110001",
"111101000101000" when"101011110010",
"111101000101010" when"101011110011",
"111101000101011" when"101011110100",
"111101000101100" when"101011110101",
"111101000101110" when"101011110110",
"111101000101111" when"101011110111",
"111101000110001" when"101011111000",
"111101000110010" when"101011111001",
"111101000110011" when"101011111010",
"111101000110101" when"101011111011",
"111101000110110" when"101011111100",
"111101000111000" when"101011111101",
"111101000111001" when"101011111110",
"111101000111010" when"101011111111",
"111101000111100" when"101100000000",
"111101000111101" when"101100000001",
"111101000111111" when"101100000010",
"111101001000000" when"101100000011",
"111101001000001" when"101100000100",
"111101001000011" when"101100000101",
"111101001000100" when"101100000110",
"111101001000110" when"101100000111",
"111101001000111" when"101100001000",
"111101001001000" when"101100001001",
"111101001001010" when"101100001010",
"111101001001011" when"101100001011",
"111101001001101" when"101100001100",
"111101001001110" when"101100001101",
"111101001001111" when"101100001110",
"111101001010001" when"101100001111",
"111101001010010" when"101100010000",
"111101001010100" when"101100010001",
"111101001010101" when"101100010010",
"111101001010110" when"101100010011",
"111101001011000" when"101100010100",
"111101001011001" when"101100010101",
"111101001011011" when"101100010110",
"111101001011100" when"101100010111",
"111101001011101" when"101100011000",
"111101001011111" when"101100011001",
"111101001100000" when"101100011010",
"111101001100001" when"101100011011",
"111101001100011" when"101100011100",
"111101001100100" when"101100011101",
"111101001100110" when"101100011110",
"111101001100111" when"101100011111",
"111101001101000" when"101100100000",
"111101001101010" when"101100100001",
"111101001101011" when"101100100010",
"111101001101101" when"101100100011",
"111101001101110" when"101100100100",
"111101001101111" when"101100100101",
"111101001110001" when"101100100110",
"111101001110010" when"101100100111",
"111101001110011" when"101100101000",
"111101001110101" when"101100101001",
"111101001110110" when"101100101010",
"111101001111000" when"101100101011",
"111101001111001" when"101100101100",
"111101001111010" when"101100101101",
"111101001111100" when"101100101110",
"111101001111101" when"101100101111",
"111101001111110" when"101100110000",
"111101010000000" when"101100110001",
"111101010000001" when"101100110010",
"111101010000011" when"101100110011",
"111101010000100" when"101100110100",
"111101010000101" when"101100110101",
"111101010000111" when"101100110110",
"111101010001000" when"101100110111",
"111101010001001" when"101100111000",
"111101010001011" when"101100111001",
"111101010001100" when"101100111010",
"111101010001110" when"101100111011",
"111101010001111" when"101100111100",
"111101010010000" when"101100111101",
"111101010010010" when"101100111110",
"111101010010011" when"101100111111",
"111101010010100" when"101101000000",
"111101010010110" when"101101000001",
"111101010010111" when"101101000010",
"111101010011000" when"101101000011",
"111101010011010" when"101101000100",
"111101010011011" when"101101000101",
"111101010011101" when"101101000110",
"111101010011110" when"101101000111",
"111101010011111" when"101101001000",
"111101010100001" when"101101001001",
"111101010100010" when"101101001010",
"111101010100011" when"101101001011",
"111101010100101" when"101101001100",
"111101010100110" when"101101001101",
"111101010100111" when"101101001110",
"111101010101001" when"101101001111",
"111101010101010" when"101101010000",
"111101010101100" when"101101010001",
"111101010101101" when"101101010010",
"111101010101110" when"101101010011",
"111101010110000" when"101101010100",
"111101010110001" when"101101010101",
"111101010110010" when"101101010110",
"111101010110100" when"101101010111",
"111101010110101" when"101101011000",
"111101010110110" when"101101011001",
"111101010111000" when"101101011010",
"111101010111001" when"101101011011",
"111101010111010" when"101101011100",
"111101010111100" when"101101011101",
"111101010111101" when"101101011110",
"111101010111111" when"101101011111",
"111101011000000" when"101101100000",
"111101011000001" when"101101100001",
"111101011000011" when"101101100010",
"111101011000100" when"101101100011",
"111101011000101" when"101101100100",
"111101011000111" when"101101100101",
"111101011001000" when"101101100110",
"111101011001001" when"101101100111",
"111101011001011" when"101101101000",
"111101011001100" when"101101101001",
"111101011001101" when"101101101010",
"111101011001111" when"101101101011",
"111101011010000" when"101101101100",
"111101011010001" when"101101101101",
"111101011010011" when"101101101110",
"111101011010100" when"101101101111",
"111101011010110" when"101101110000",
"111101011010111" when"101101110001",
"111101011011000" when"101101110010",
"111101011011010" when"101101110011",
"111101011011011" when"101101110100",
"111101011011100" when"101101110101",
"111101011011110" when"101101110110",
"111101011011111" when"101101110111",
"111101011100000" when"101101111000",
"111101011100010" when"101101111001",
"111101011100011" when"101101111010",
"111101011100100" when"101101111011",
"111101011100110" when"101101111100",
"111101011100111" when"101101111101",
"111101011101000" when"101101111110",
"111101011101010" when"101101111111",
"111101011101011" when"101110000000",
"111101011101100" when"101110000001",
"111101011101110" when"101110000010",
"111101011101111" when"101110000011",
"111101011110000" when"101110000100",
"111101011110010" when"101110000101",
"111101011110011" when"101110000110",
"111101011110100" when"101110000111",
"111101011110110" when"101110001000",
"111101011110111" when"101110001001",
"111101011111000" when"101110001010",
"111101011111010" when"101110001011",
"111101011111011" when"101110001100",
"111101011111100" when"101110001101",
"111101011111110" when"101110001110",
"111101011111111" when"101110001111",
"111101100000000" when"101110010000",
"111101100000010" when"101110010001",
"111101100000011" when"101110010010",
"111101100000100" when"101110010011",
"111101100000110" when"101110010100",
"111101100000111" when"101110010101",
"111101100001000" when"101110010110",
"111101100001010" when"101110010111",
"111101100001011" when"101110011000",
"111101100001100" when"101110011001",
"111101100001110" when"101110011010",
"111101100001111" when"101110011011",
"111101100010000" when"101110011100",
"111101100010010" when"101110011101",
"111101100010011" when"101110011110",
"111101100010100" when"101110011111",
"111101100010110" when"101110100000",
"111101100010111" when"101110100001",
"111101100011000" when"101110100010",
"111101100011010" when"101110100011",
"111101100011011" when"101110100100",
"111101100011100" when"101110100101",
"111101100011101" when"101110100110",
"111101100011111" when"101110100111",
"111101100100000" when"101110101000",
"111101100100001" when"101110101001",
"111101100100011" when"101110101010",
"111101100100100" when"101110101011",
"111101100100101" when"101110101100",
"111101100100111" when"101110101101",
"111101100101000" when"101110101110",
"111101100101001" when"101110101111",
"111101100101011" when"101110110000",
"111101100101100" when"101110110001",
"111101100101101" when"101110110010",
"111101100101111" when"101110110011",
"111101100110000" when"101110110100",
"111101100110001" when"101110110101",
"111101100110011" when"101110110110",
"111101100110100" when"101110110111",
"111101100110101" when"101110111000",
"111101100110111" when"101110111001",
"111101100111000" when"101110111010",
"111101100111001" when"101110111011",
"111101100111010" when"101110111100",
"111101100111100" when"101110111101",
"111101100111101" when"101110111110",
"111101100111110" when"101110111111",
"111101101000000" when"101111000000",
"111101101000001" when"101111000001",
"111101101000010" when"101111000010",
"111101101000100" when"101111000011",
"111101101000101" when"101111000100",
"111101101000110" when"101111000101",
"111101101001000" when"101111000110",
"111101101001001" when"101111000111",
"111101101001010" when"101111001000",
"111101101001011" when"101111001001",
"111101101001101" when"101111001010",
"111101101001110" when"101111001011",
"111101101001111" when"101111001100",
"111101101010001" when"101111001101",
"111101101010010" when"101111001110",
"111101101010011" when"101111001111",
"111101101010101" when"101111010000",
"111101101010110" when"101111010001",
"111101101010111" when"101111010010",
"111101101011000" when"101111010011",
"111101101011010" when"101111010100",
"111101101011011" when"101111010101",
"111101101011100" when"101111010110",
"111101101011110" when"101111010111",
"111101101011111" when"101111011000",
"111101101100000" when"101111011001",
"111101101100010" when"101111011010",
"111101101100011" when"101111011011",
"111101101100100" when"101111011100",
"111101101100101" when"101111011101",
"111101101100111" when"101111011110",
"111101101101000" when"101111011111",
"111101101101001" when"101111100000",
"111101101101011" when"101111100001",
"111101101101100" when"101111100010",
"111101101101101" when"101111100011",
"111101101101111" when"101111100100",
"111101101110000" when"101111100101",
"111101101110001" when"101111100110",
"111101101110010" when"101111100111",
"111101101110100" when"101111101000",
"111101101110101" when"101111101001",
"111101101110110" when"101111101010",
"111101101111000" when"101111101011",
"111101101111001" when"101111101100",
"111101101111010" when"101111101101",
"111101101111011" when"101111101110",
"111101101111101" when"101111101111",
"111101101111110" when"101111110000",
"111101101111111" when"101111110001",
"111101110000001" when"101111110010",
"111101110000010" when"101111110011",
"111101110000011" when"101111110100",
"111101110000101" when"101111110101",
"111101110000110" when"101111110110",
"111101110000111" when"101111110111",
"111101110001000" when"101111111000",
"111101110001010" when"101111111001",
"111101110001011" when"101111111010",
"111101110001100" when"101111111011",
"111101110001110" when"101111111100",
"111101110001111" when"101111111101",
"111101110010000" when"101111111110",
"111101110010001" when"101111111111",
"111101110010011" when"110000000000",
"111101110010100" when"110000000001",
"111101110010101" when"110000000010",
"111101110010110" when"110000000011",
"111101110011000" when"110000000100",
"111101110011001" when"110000000101",
"111101110011010" when"110000000110",
"111101110011100" when"110000000111",
"111101110011101" when"110000001000",
"111101110011110" when"110000001001",
"111101110011111" when"110000001010",
"111101110100001" when"110000001011",
"111101110100010" when"110000001100",
"111101110100011" when"110000001101",
"111101110100101" when"110000001110",
"111101110100110" when"110000001111",
"111101110100111" when"110000010000",
"111101110101000" when"110000010001",
"111101110101010" when"110000010010",
"111101110101011" when"110000010011",
"111101110101100" when"110000010100",
"111101110101101" when"110000010101",
"111101110101111" when"110000010110",
"111101110110000" when"110000010111",
"111101110110001" when"110000011000",
"111101110110011" when"110000011001",
"111101110110100" when"110000011010",
"111101110110101" when"110000011011",
"111101110110110" when"110000011100",
"111101110111000" when"110000011101",
"111101110111001" when"110000011110",
"111101110111010" when"110000011111",
"111101110111011" when"110000100000",
"111101110111101" when"110000100001",
"111101110111110" when"110000100010",
"111101110111111" when"110000100011",
"111101111000001" when"110000100100",
"111101111000010" when"110000100101",
"111101111000011" when"110000100110",
"111101111000100" when"110000100111",
"111101111000110" when"110000101000",
"111101111000111" when"110000101001",
"111101111001000" when"110000101010",
"111101111001001" when"110000101011",
"111101111001011" when"110000101100",
"111101111001100" when"110000101101",
"111101111001101" when"110000101110",
"111101111001110" when"110000101111",
"111101111010000" when"110000110000",
"111101111010001" when"110000110001",
"111101111010010" when"110000110010",
"111101111010011" when"110000110011",
"111101111010101" when"110000110100",
"111101111010110" when"110000110101",
"111101111010111" when"110000110110",
"111101111011001" when"110000110111",
"111101111011010" when"110000111000",
"111101111011011" when"110000111001",
"111101111011100" when"110000111010",
"111101111011110" when"110000111011",
"111101111011111" when"110000111100",
"111101111100000" when"110000111101",
"111101111100001" when"110000111110",
"111101111100011" when"110000111111",
"111101111100100" when"110001000000",
"111101111100101" when"110001000001",
"111101111100110" when"110001000010",
"111101111101000" when"110001000011",
"111101111101001" when"110001000100",
"111101111101010" when"110001000101",
"111101111101011" when"110001000110",
"111101111101101" when"110001000111",
"111101111101110" when"110001001000",
"111101111101111" when"110001001001",
"111101111110000" when"110001001010",
"111101111110010" when"110001001011",
"111101111110011" when"110001001100",
"111101111110100" when"110001001101",
"111101111110101" when"110001001110",
"111101111110111" when"110001001111",
"111101111111000" when"110001010000",
"111101111111001" when"110001010001",
"111101111111010" when"110001010010",
"111101111111100" when"110001010011",
"111101111111101" when"110001010100",
"111101111111110" when"110001010101",
"111101111111111" when"110001010110",
"111110000000001" when"110001010111",
"111110000000010" when"110001011000",
"111110000000011" when"110001011001",
"111110000000100" when"110001011010",
"111110000000110" when"110001011011",
"111110000000111" when"110001011100",
"111110000001000" when"110001011101",
"111110000001001" when"110001011110",
"111110000001011" when"110001011111",
"111110000001100" when"110001100000",
"111110000001101" when"110001100001",
"111110000001110" when"110001100010",
"111110000010000" when"110001100011",
"111110000010001" when"110001100100",
"111110000010010" when"110001100101",
"111110000010011" when"110001100110",
"111110000010101" when"110001100111",
"111110000010110" when"110001101000",
"111110000010111" when"110001101001",
"111110000011000" when"110001101010",
"111110000011010" when"110001101011",
"111110000011011" when"110001101100",
"111110000011100" when"110001101101",
"111110000011101" when"110001101110",
"111110000011110" when"110001101111",
"111110000100000" when"110001110000",
"111110000100001" when"110001110001",
"111110000100010" when"110001110010",
"111110000100011" when"110001110011",
"111110000100101" when"110001110100",
"111110000100110" when"110001110101",
"111110000100111" when"110001110110",
"111110000101000" when"110001110111",
"111110000101010" when"110001111000",
"111110000101011" when"110001111001",
"111110000101100" when"110001111010",
"111110000101101" when"110001111011",
"111110000101111" when"110001111100",
"111110000110000" when"110001111101",
"111110000110001" when"110001111110",
"111110000110010" when"110001111111",
"111110000110011" when"110010000000",
"111110000110101" when"110010000001",
"111110000110110" when"110010000010",
"111110000110111" when"110010000011",
"111110000111000" when"110010000100",
"111110000111010" when"110010000101",
"111110000111011" when"110010000110",
"111110000111100" when"110010000111",
"111110000111101" when"110010001000",
"111110000111111" when"110010001001",
"111110001000000" when"110010001010",
"111110001000001" when"110010001011",
"111110001000010" when"110010001100",
"111110001000011" when"110010001101",
"111110001000101" when"110010001110",
"111110001000110" when"110010001111",
"111110001000111" when"110010010000",
"111110001001000" when"110010010001",
"111110001001010" when"110010010010",
"111110001001011" when"110010010011",
"111110001001100" when"110010010100",
"111110001001101" when"110010010101",
"111110001001110" when"110010010110",
"111110001010000" when"110010010111",
"111110001010001" when"110010011000",
"111110001010010" when"110010011001",
"111110001010011" when"110010011010",
"111110001010101" when"110010011011",
"111110001010110" when"110010011100",
"111110001010111" when"110010011101",
"111110001011000" when"110010011110",
"111110001011001" when"110010011111",
"111110001011011" when"110010100000",
"111110001011100" when"110010100001",
"111110001011101" when"110010100010",
"111110001011110" when"110010100011",
"111110001100000" when"110010100100",
"111110001100001" when"110010100101",
"111110001100010" when"110010100110",
"111110001100011" when"110010100111",
"111110001100100" when"110010101000",
"111110001100110" when"110010101001",
"111110001100111" when"110010101010",
"111110001101000" when"110010101011",
"111110001101001" when"110010101100",
"111110001101010" when"110010101101",
"111110001101100" when"110010101110",
"111110001101101" when"110010101111",
"111110001101110" when"110010110000",
"111110001101111" when"110010110001",
"111110001110001" when"110010110010",
"111110001110010" when"110010110011",
"111110001110011" when"110010110100",
"111110001110100" when"110010110101",
"111110001110101" when"110010110110",
"111110001110111" when"110010110111",
"111110001111000" when"110010111000",
"111110001111001" when"110010111001",
"111110001111010" when"110010111010",
"111110001111011" when"110010111011",
"111110001111101" when"110010111100",
"111110001111110" when"110010111101",
"111110001111111" when"110010111110",
"111110010000000" when"110010111111",
"111110010000001" when"110011000000",
"111110010000011" when"110011000001",
"111110010000100" when"110011000010",
"111110010000101" when"110011000011",
"111110010000110" when"110011000100",
"111110010000111" when"110011000101",
"111110010001001" when"110011000110",
"111110010001010" when"110011000111",
"111110010001011" when"110011001000",
"111110010001100" when"110011001001",
"111110010001110" when"110011001010",
"111110010001111" when"110011001011",
"111110010010000" when"110011001100",
"111110010010001" when"110011001101",
"111110010010010" when"110011001110",
"111110010010100" when"110011001111",
"111110010010101" when"110011010000",
"111110010010110" when"110011010001",
"111110010010111" when"110011010010",
"111110010011000" when"110011010011",
"111110010011010" when"110011010100",
"111110010011011" when"110011010101",
"111110010011100" when"110011010110",
"111110010011101" when"110011010111",
"111110010011110" when"110011011000",
"111110010100000" when"110011011001",
"111110010100001" when"110011011010",
"111110010100010" when"110011011011",
"111110010100011" when"110011011100",
"111110010100100" when"110011011101",
"111110010100110" when"110011011110",
"111110010100111" when"110011011111",
"111110010101000" when"110011100000",
"111110010101001" when"110011100001",
"111110010101010" when"110011100010",
"111110010101011" when"110011100011",
"111110010101101" when"110011100100",
"111110010101110" when"110011100101",
"111110010101111" when"110011100110",
"111110010110000" when"110011100111",
"111110010110001" when"110011101000",
"111110010110011" when"110011101001",
"111110010110100" when"110011101010",
"111110010110101" when"110011101011",
"111110010110110" when"110011101100",
"111110010110111" when"110011101101",
"111110010111001" when"110011101110",
"111110010111010" when"110011101111",
"111110010111011" when"110011110000",
"111110010111100" when"110011110001",
"111110010111101" when"110011110010",
"111110010111111" when"110011110011",
"111110011000000" when"110011110100",
"111110011000001" when"110011110101",
"111110011000010" when"110011110110",
"111110011000011" when"110011110111",
"111110011000100" when"110011111000",
"111110011000110" when"110011111001",
"111110011000111" when"110011111010",
"111110011001000" when"110011111011",
"111110011001001" when"110011111100",
"111110011001010" when"110011111101",
"111110011001100" when"110011111110",
"111110011001101" when"110011111111",
"111110011001110" when"110100000000",
"111110011001111" when"110100000001",
"111110011010000" when"110100000010",
"111110011010010" when"110100000011",
"111110011010011" when"110100000100",
"111110011010100" when"110100000101",
"111110011010101" when"110100000110",
"111110011010110" when"110100000111",
"111110011010111" when"110100001000",
"111110011011001" when"110100001001",
"111110011011010" when"110100001010",
"111110011011011" when"110100001011",
"111110011011100" when"110100001100",
"111110011011101" when"110100001101",
"111110011011111" when"110100001110",
"111110011100000" when"110100001111",
"111110011100001" when"110100010000",
"111110011100010" when"110100010001",
"111110011100011" when"110100010010",
"111110011100100" when"110100010011",
"111110011100110" when"110100010100",
"111110011100111" when"110100010101",
"111110011101000" when"110100010110",
"111110011101001" when"110100010111",
"111110011101010" when"110100011000",
"111110011101011" when"110100011001",
"111110011101101" when"110100011010",
"111110011101110" when"110100011011",
"111110011101111" when"110100011100",
"111110011110000" when"110100011101",
"111110011110001" when"110100011110",
"111110011110010" when"110100011111",
"111110011110100" when"110100100000",
"111110011110101" when"110100100001",
"111110011110110" when"110100100010",
"111110011110111" when"110100100011",
"111110011111000" when"110100100100",
"111110011111010" when"110100100101",
"111110011111011" when"110100100110",
"111110011111100" when"110100100111",
"111110011111101" when"110100101000",
"111110011111110" when"110100101001",
"111110011111111" when"110100101010",
"111110100000001" when"110100101011",
"111110100000010" when"110100101100",
"111110100000011" when"110100101101",
"111110100000100" when"110100101110",
"111110100000101" when"110100101111",
"111110100000110" when"110100110000",
"111110100001000" when"110100110001",
"111110100001001" when"110100110010",
"111110100001010" when"110100110011",
"111110100001011" when"110100110100",
"111110100001100" when"110100110101",
"111110100001101" when"110100110110",
"111110100001111" when"110100110111",
"111110100010000" when"110100111000",
"111110100010001" when"110100111001",
"111110100010010" when"110100111010",
"111110100010011" when"110100111011",
"111110100010100" when"110100111100",
"111110100010110" when"110100111101",
"111110100010111" when"110100111110",
"111110100011000" when"110100111111",
"111110100011001" when"110101000000",
"111110100011010" when"110101000001",
"111110100011011" when"110101000010",
"111110100011100" when"110101000011",
"111110100011110" when"110101000100",
"111110100011111" when"110101000101",
"111110100100000" when"110101000110",
"111110100100001" when"110101000111",
"111110100100010" when"110101001000",
"111110100100011" when"110101001001",
"111110100100101" when"110101001010",
"111110100100110" when"110101001011",
"111110100100111" when"110101001100",
"111110100101000" when"110101001101",
"111110100101001" when"110101001110",
"111110100101010" when"110101001111",
"111110100101100" when"110101010000",
"111110100101101" when"110101010001",
"111110100101110" when"110101010010",
"111110100101111" when"110101010011",
"111110100110000" when"110101010100",
"111110100110001" when"110101010101",
"111110100110010" when"110101010110",
"111110100110100" when"110101010111",
"111110100110101" when"110101011000",
"111110100110110" when"110101011001",
"111110100110111" when"110101011010",
"111110100111000" when"110101011011",
"111110100111001" when"110101011100",
"111110100111011" when"110101011101",
"111110100111100" when"110101011110",
"111110100111101" when"110101011111",
"111110100111110" when"110101100000",
"111110100111111" when"110101100001",
"111110101000000" when"110101100010",
"111110101000001" when"110101100011",
"111110101000011" when"110101100100",
"111110101000100" when"110101100101",
"111110101000101" when"110101100110",
"111110101000110" when"110101100111",
"111110101000111" when"110101101000",
"111110101001000" when"110101101001",
"111110101001001" when"110101101010",
"111110101001011" when"110101101011",
"111110101001100" when"110101101100",
"111110101001101" when"110101101101",
"111110101001110" when"110101101110",
"111110101001111" when"110101101111",
"111110101010000" when"110101110000",
"111110101010010" when"110101110001",
"111110101010011" when"110101110010",
"111110101010100" when"110101110011",
"111110101010101" when"110101110100",
"111110101010110" when"110101110101",
"111110101010111" when"110101110110",
"111110101011000" when"110101110111",
"111110101011010" when"110101111000",
"111110101011011" when"110101111001",
"111110101011100" when"110101111010",
"111110101011101" when"110101111011",
"111110101011110" when"110101111100",
"111110101011111" when"110101111101",
"111110101100000" when"110101111110",
"111110101100010" when"110101111111",
"111110101100011" when"110110000000",
"111110101100100" when"110110000001",
"111110101100101" when"110110000010",
"111110101100110" when"110110000011",
"111110101100111" when"110110000100",
"111110101101000" when"110110000101",
"111110101101001" when"110110000110",
"111110101101011" when"110110000111",
"111110101101100" when"110110001000",
"111110101101101" when"110110001001",
"111110101101110" when"110110001010",
"111110101101111" when"110110001011",
"111110101110000" when"110110001100",
"111110101110001" when"110110001101",
"111110101110011" when"110110001110",
"111110101110100" when"110110001111",
"111110101110101" when"110110010000",
"111110101110110" when"110110010001",
"111110101110111" when"110110010010",
"111110101111000" when"110110010011",
"111110101111001" when"110110010100",
"111110101111011" when"110110010101",
"111110101111100" when"110110010110",
"111110101111101" when"110110010111",
"111110101111110" when"110110011000",
"111110101111111" when"110110011001",
"111110110000000" when"110110011010",
"111110110000001" when"110110011011",
"111110110000010" when"110110011100",
"111110110000100" when"110110011101",
"111110110000101" when"110110011110",
"111110110000110" when"110110011111",
"111110110000111" when"110110100000",
"111110110001000" when"110110100001",
"111110110001001" when"110110100010",
"111110110001010" when"110110100011",
"111110110001011" when"110110100100",
"111110110001101" when"110110100101",
"111110110001110" when"110110100110",
"111110110001111" when"110110100111",
"111110110010000" when"110110101000",
"111110110010001" when"110110101001",
"111110110010010" when"110110101010",
"111110110010011" when"110110101011",
"111110110010100" when"110110101100",
"111110110010110" when"110110101101",
"111110110010111" when"110110101110",
"111110110011000" when"110110101111",
"111110110011001" when"110110110000",
"111110110011010" when"110110110001",
"111110110011011" when"110110110010",
"111110110011100" when"110110110011",
"111110110011101" when"110110110100",
"111110110011111" when"110110110101",
"111110110100000" when"110110110110",
"111110110100001" when"110110110111",
"111110110100010" when"110110111000",
"111110110100011" when"110110111001",
"111110110100100" when"110110111010",
"111110110100101" when"110110111011",
"111110110100110" when"110110111100",
"111110110101000" when"110110111101",
"111110110101001" when"110110111110",
"111110110101010" when"110110111111",
"111110110101011" when"110111000000",
"111110110101100" when"110111000001",
"111110110101101" when"110111000010",
"111110110101110" when"110111000011",
"111110110101111" when"110111000100",
"111110110110001" when"110111000101",
"111110110110010" when"110111000110",
"111110110110011" when"110111000111",
"111110110110100" when"110111001000",
"111110110110101" when"110111001001",
"111110110110110" when"110111001010",
"111110110110111" when"110111001011",
"111110110111000" when"110111001100",
"111110110111001" when"110111001101",
"111110110111011" when"110111001110",
"111110110111100" when"110111001111",
"111110110111101" when"110111010000",
"111110110111110" when"110111010001",
"111110110111111" when"110111010010",
"111110111000000" when"110111010011",
"111110111000001" when"110111010100",
"111110111000010" when"110111010101",
"111110111000011" when"110111010110",
"111110111000101" when"110111010111",
"111110111000110" when"110111011000",
"111110111000111" when"110111011001",
"111110111001000" when"110111011010",
"111110111001001" when"110111011011",
"111110111001010" when"110111011100",
"111110111001011" when"110111011101",
"111110111001100" when"110111011110",
"111110111001101" when"110111011111",
"111110111001111" when"110111100000",
"111110111010000" when"110111100001",
"111110111010001" when"110111100010",
"111110111010010" when"110111100011",
"111110111010011" when"110111100100",
"111110111010100" when"110111100101",
"111110111010101" when"110111100110",
"111110111010110" when"110111100111",
"111110111010111" when"110111101000",
"111110111011001" when"110111101001",
"111110111011010" when"110111101010",
"111110111011011" when"110111101011",
"111110111011100" when"110111101100",
"111110111011101" when"110111101101",
"111110111011110" when"110111101110",
"111110111011111" when"110111101111",
"111110111100000" when"110111110000",
"111110111100001" when"110111110001",
"111110111100010" when"110111110010",
"111110111100100" when"110111110011",
"111110111100101" when"110111110100",
"111110111100110" when"110111110101",
"111110111100111" when"110111110110",
"111110111101000" when"110111110111",
"111110111101001" when"110111111000",
"111110111101010" when"110111111001",
"111110111101011" when"110111111010",
"111110111101100" when"110111111011",
"111110111101110" when"110111111100",
"111110111101111" when"110111111101",
"111110111110000" when"110111111110",
"111110111110001" when"110111111111",
"111110111110010" when"111000000000",
"111110111110011" when"111000000001",
"111110111110100" when"111000000010",
"111110111110101" when"111000000011",
"111110111110110" when"111000000100",
"111110111110111" when"111000000101",
"111110111111001" when"111000000110",
"111110111111010" when"111000000111",
"111110111111011" when"111000001000",
"111110111111100" when"111000001001",
"111110111111101" when"111000001010",
"111110111111110" when"111000001011",
"111110111111111" when"111000001100",
"111111000000000" when"111000001101",
"111111000000001" when"111000001110",
"111111000000010" when"111000001111",
"111111000000011" when"111000010000",
"111111000000101" when"111000010001",
"111111000000110" when"111000010010",
"111111000000111" when"111000010011",
"111111000001000" when"111000010100",
"111111000001001" when"111000010101",
"111111000001010" when"111000010110",
"111111000001011" when"111000010111",
"111111000001100" when"111000011000",
"111111000001101" when"111000011001",
"111111000001110" when"111000011010",
"111111000001111" when"111000011011",
"111111000010001" when"111000011100",
"111111000010010" when"111000011101",
"111111000010011" when"111000011110",
"111111000010100" when"111000011111",
"111111000010101" when"111000100000",
"111111000010110" when"111000100001",
"111111000010111" when"111000100010",
"111111000011000" when"111000100011",
"111111000011001" when"111000100100",
"111111000011010" when"111000100101",
"111111000011011" when"111000100110",
"111111000011101" when"111000100111",
"111111000011110" when"111000101000",
"111111000011111" when"111000101001",
"111111000100000" when"111000101010",
"111111000100001" when"111000101011",
"111111000100010" when"111000101100",
"111111000100011" when"111000101101",
"111111000100100" when"111000101110",
"111111000100101" when"111000101111",
"111111000100110" when"111000110000",
"111111000100111" when"111000110001",
"111111000101000" when"111000110010",
"111111000101010" when"111000110011",
"111111000101011" when"111000110100",
"111111000101100" when"111000110101",
"111111000101101" when"111000110110",
"111111000101110" when"111000110111",
"111111000101111" when"111000111000",
"111111000110000" when"111000111001",
"111111000110001" when"111000111010",
"111111000110010" when"111000111011",
"111111000110011" when"111000111100",
"111111000110100" when"111000111101",
"111111000110101" when"111000111110",
"111111000110111" when"111000111111",
"111111000111000" when"111001000000",
"111111000111001" when"111001000001",
"111111000111010" when"111001000010",
"111111000111011" when"111001000011",
"111111000111100" when"111001000100",
"111111000111101" when"111001000101",
"111111000111110" when"111001000110",
"111111000111111" when"111001000111",
"111111001000000" when"111001001000",
"111111001000001" when"111001001001",
"111111001000010" when"111001001010",
"111111001000100" when"111001001011",
"111111001000101" when"111001001100",
"111111001000110" when"111001001101",
"111111001000111" when"111001001110",
"111111001001000" when"111001001111",
"111111001001001" when"111001010000",
"111111001001010" when"111001010001",
"111111001001011" when"111001010010",
"111111001001100" when"111001010011",
"111111001001101" when"111001010100",
"111111001001110" when"111001010101",
"111111001001111" when"111001010110",
"111111001010000" when"111001010111",
"111111001010001" when"111001011000",
"111111001010011" when"111001011001",
"111111001010100" when"111001011010",
"111111001010101" when"111001011011",
"111111001010110" when"111001011100",
"111111001010111" when"111001011101",
"111111001011000" when"111001011110",
"111111001011001" when"111001011111",
"111111001011010" when"111001100000",
"111111001011011" when"111001100001",
"111111001011100" when"111001100010",
"111111001011101" when"111001100011",
"111111001011110" when"111001100100",
"111111001011111" when"111001100101",
"111111001100000" when"111001100110",
"111111001100010" when"111001100111",
"111111001100011" when"111001101000",
"111111001100100" when"111001101001",
"111111001100101" when"111001101010",
"111111001100110" when"111001101011",
"111111001100111" when"111001101100",
"111111001101000" when"111001101101",
"111111001101001" when"111001101110",
"111111001101010" when"111001101111",
"111111001101011" when"111001110000",
"111111001101100" when"111001110001",
"111111001101101" when"111001110010",
"111111001101110" when"111001110011",
"111111001101111" when"111001110100",
"111111001110000" when"111001110101",
"111111001110010" when"111001110110",
"111111001110011" when"111001110111",
"111111001110100" when"111001111000",
"111111001110101" when"111001111001",
"111111001110110" when"111001111010",
"111111001110111" when"111001111011",
"111111001111000" when"111001111100",
"111111001111001" when"111001111101",
"111111001111010" when"111001111110",
"111111001111011" when"111001111111",
"111111001111100" when"111010000000",
"111111001111101" when"111010000001",
"111111001111110" when"111010000010",
"111111001111111" when"111010000011",
"111111010000000" when"111010000100",
"111111010000001" when"111010000101",
"111111010000011" when"111010000110",
"111111010000100" when"111010000111",
"111111010000101" when"111010001000",
"111111010000110" when"111010001001",
"111111010000111" when"111010001010",
"111111010001000" when"111010001011",
"111111010001001" when"111010001100",
"111111010001010" when"111010001101",
"111111010001011" when"111010001110",
"111111010001100" when"111010001111",
"111111010001101" when"111010010000",
"111111010001110" when"111010010001",
"111111010001111" when"111010010010",
"111111010010000" when"111010010011",
"111111010010001" when"111010010100",
"111111010010010" when"111010010101",
"111111010010011" when"111010010110",
"111111010010100" when"111010010111",
"111111010010110" when"111010011000",
"111111010010111" when"111010011001",
"111111010011000" when"111010011010",
"111111010011001" when"111010011011",
"111111010011010" when"111010011100",
"111111010011011" when"111010011101",
"111111010011100" when"111010011110",
"111111010011101" when"111010011111",
"111111010011110" when"111010100000",
"111111010011111" when"111010100001",
"111111010100000" when"111010100010",
"111111010100001" when"111010100011",
"111111010100010" when"111010100100",
"111111010100011" when"111010100101",
"111111010100100" when"111010100110",
"111111010100101" when"111010100111",
"111111010100110" when"111010101000",
"111111010100111" when"111010101001",
"111111010101000" when"111010101010",
"111111010101010" when"111010101011",
"111111010101011" when"111010101100",
"111111010101100" when"111010101101",
"111111010101101" when"111010101110",
"111111010101110" when"111010101111",
"111111010101111" when"111010110000",
"111111010110000" when"111010110001",
"111111010110001" when"111010110010",
"111111010110010" when"111010110011",
"111111010110011" when"111010110100",
"111111010110100" when"111010110101",
"111111010110101" when"111010110110",
"111111010110110" when"111010110111",
"111111010110111" when"111010111000",
"111111010111000" when"111010111001",
"111111010111001" when"111010111010",
"111111010111010" when"111010111011",
"111111010111011" when"111010111100",
"111111010111100" when"111010111101",
"111111010111101" when"111010111110",
"111111010111110" when"111010111111",
"111111010111111" when"111011000000",
"111111011000001" when"111011000001",
"111111011000010" when"111011000010",
"111111011000011" when"111011000011",
"111111011000100" when"111011000100",
"111111011000101" when"111011000101",
"111111011000110" when"111011000110",
"111111011000111" when"111011000111",
"111111011001000" when"111011001000",
"111111011001001" when"111011001001",
"111111011001010" when"111011001010",
"111111011001011" when"111011001011",
"111111011001100" when"111011001100",
"111111011001101" when"111011001101",
"111111011001110" when"111011001110",
"111111011001111" when"111011001111",
"111111011010000" when"111011010000",
"111111011010001" when"111011010001",
"111111011010010" when"111011010010",
"111111011010011" when"111011010011",
"111111011010100" when"111011010100",
"111111011010101" when"111011010101",
"111111011010110" when"111011010110",
"111111011010111" when"111011010111",
"111111011011000" when"111011011000",
"111111011011001" when"111011011001",
"111111011011011" when"111011011010",
"111111011011100" when"111011011011",
"111111011011101" when"111011011100",
"111111011011110" when"111011011101",
"111111011011111" when"111011011110",
"111111011100000" when"111011011111",
"111111011100001" when"111011100000",
"111111011100010" when"111011100001",
"111111011100011" when"111011100010",
"111111011100100" when"111011100011",
"111111011100101" when"111011100100",
"111111011100110" when"111011100101",
"111111011100111" when"111011100110",
"111111011101000" when"111011100111",
"111111011101001" when"111011101000",
"111111011101010" when"111011101001",
"111111011101011" when"111011101010",
"111111011101100" when"111011101011",
"111111011101101" when"111011101100",
"111111011101110" when"111011101101",
"111111011101111" when"111011101110",
"111111011110000" when"111011101111",
"111111011110001" when"111011110000",
"111111011110010" when"111011110001",
"111111011110011" when"111011110010",
"111111011110100" when"111011110011",
"111111011110101" when"111011110100",
"111111011110110" when"111011110101",
"111111011110111" when"111011110110",
"111111011111000" when"111011110111",
"111111011111001" when"111011111000",
"111111011111011" when"111011111001",
"111111011111100" when"111011111010",
"111111011111101" when"111011111011",
"111111011111110" when"111011111100",
"111111011111111" when"111011111101",
"111111100000000" when"111011111110",
"111111100000001" when"111011111111",
"111111100000010" when"111100000000",
"111111100000011" when"111100000001",
"111111100000100" when"111100000010",
"111111100000101" when"111100000011",
"111111100000110" when"111100000100",
"111111100000111" when"111100000101",
"111111100001000" when"111100000110",
"111111100001001" when"111100000111",
"111111100001010" when"111100001000",
"111111100001011" when"111100001001",
"111111100001100" when"111100001010",
"111111100001101" when"111100001011",
"111111100001110" when"111100001100",
"111111100001111" when"111100001101",
"111111100010000" when"111100001110",
"111111100010001" when"111100001111",
"111111100010010" when"111100010000",
"111111100010011" when"111100010001",
"111111100010100" when"111100010010",
"111111100010101" when"111100010011",
"111111100010110" when"111100010100",
"111111100010111" when"111100010101",
"111111100011000" when"111100010110",
"111111100011001" when"111100010111",
"111111100011010" when"111100011000",
"111111100011011" when"111100011001",
"111111100011100" when"111100011010",
"111111100011101" when"111100011011",
"111111100011110" when"111100011100",
"111111100011111" when"111100011101",
"111111100100000" when"111100011110",
"111111100100001" when"111100011111",
"111111100100010" when"111100100000",
"111111100100011" when"111100100001",
"111111100100100" when"111100100010",
"111111100100101" when"111100100011",
"111111100100110" when"111100100100",
"111111100100111" when"111100100101",
"111111100101001" when"111100100110",
"111111100101010" when"111100100111",
"111111100101011" when"111100101000",
"111111100101100" when"111100101001",
"111111100101101" when"111100101010",
"111111100101110" when"111100101011",
"111111100101111" when"111100101100",
"111111100110000" when"111100101101",
"111111100110001" when"111100101110",
"111111100110010" when"111100101111",
"111111100110011" when"111100110000",
"111111100110100" when"111100110001",
"111111100110101" when"111100110010",
"111111100110110" when"111100110011",
"111111100110111" when"111100110100",
"111111100111000" when"111100110101",
"111111100111001" when"111100110110",
"111111100111010" when"111100110111",
"111111100111011" when"111100111000",
"111111100111100" when"111100111001",
"111111100111101" when"111100111010",
"111111100111110" when"111100111011",
"111111100111111" when"111100111100",
"111111101000000" when"111100111101",
"111111101000001" when"111100111110",
"111111101000010" when"111100111111",
"111111101000011" when"111101000000",
"111111101000100" when"111101000001",
"111111101000101" when"111101000010",
"111111101000110" when"111101000011",
"111111101000111" when"111101000100",
"111111101001000" when"111101000101",
"111111101001001" when"111101000110",
"111111101001010" when"111101000111",
"111111101001011" when"111101001000",
"111111101001100" when"111101001001",
"111111101001101" when"111101001010",
"111111101001110" when"111101001011",
"111111101001111" when"111101001100",
"111111101010000" when"111101001101",
"111111101010001" when"111101001110",
"111111101010010" when"111101001111",
"111111101010011" when"111101010000",
"111111101010100" when"111101010001",
"111111101010101" when"111101010010",
"111111101010110" when"111101010011",
"111111101010111" when"111101010100",
"111111101011000" when"111101010101",
"111111101011001" when"111101010110",
"111111101011010" when"111101010111",
"111111101011011" when"111101011000",
"111111101011100" when"111101011001",
"111111101011101" when"111101011010",
"111111101011110" when"111101011011",
"111111101011111" when"111101011100",
"111111101100000" when"111101011101",
"111111101100001" when"111101011110",
"111111101100010" when"111101011111",
"111111101100011" when"111101100000",
"111111101100100" when"111101100001",
"111111101100101" when"111101100010",
"111111101100110" when"111101100011",
"111111101100111" when"111101100100",
"111111101101000" when"111101100101",
"111111101101001" when"111101100110",
"111111101101010" when"111101100111",
"111111101101011" when"111101101000",
"111111101101100" when"111101101001",
"111111101101101" when"111101101010",
"111111101101110" when"111101101011",
"111111101101111" when"111101101100",
"111111101110000" when"111101101101",
"111111101110001" when"111101101110",
"111111101110010" when"111101101111",
"111111101110011" when"111101110000",
"111111101110100" when"111101110001",
"111111101110101" when"111101110010",
"111111101110110" when"111101110011",
"111111101110111" when"111101110100",
"111111101111000" when"111101110101",
"111111101111001" when"111101110110",
"111111101111010" when"111101110111",
"111111101111011" when"111101111000",
"111111101111100" when"111101111001",
"111111101111101" when"111101111010",
"111111101111110" when"111101111011",
"111111101111111" when"111101111100",
"111111110000000" when"111101111101",
"111111110000001" when"111101111110",
"111111110000010" when"111101111111",
"111111110000011" when"111110000000",
"111111110000100" when"111110000001",
"111111110000101" when"111110000010",
"111111110000110" when"111110000011",
"111111110000111" when"111110000100",
"111111110001000" when"111110000101",
"111111110001001" when"111110000110",
"111111110001010" when"111110000111",
"111111110001011" when"111110001000",
"111111110001100" when"111110001001",
"111111110001101" when"111110001010",
"111111110001110" when"111110001011",
"111111110001111" when"111110001100",
"111111110010000" when"111110001101",
"111111110010001" when"111110001110",
"111111110010010" when"111110001111",
"111111110010011" when"111110010000",
"111111110010100" when"111110010001",
"111111110010101" when"111110010010",
"111111110010110" when"111110010011",
"111111110010111" when"111110010100",
"111111110011000" when"111110010101",
"111111110011001" when"111110010110",
"111111110011010" when"111110010111",
"111111110011011" when"111110011000",
"111111110011100" when"111110011001",
"111111110011101" when"111110011010",
"111111110011110" when"111110011011",
"111111110011111" when"111110011100",
"111111110100000" when"111110011101",
"111111110100001" when"111110011110",
"111111110100010" when"111110011111",
"111111110100011" when"111110100000",
"111111110100100" when"111110100001",
"111111110100100" when"111110100010",
"111111110100101" when"111110100011",
"111111110100110" when"111110100100",
"111111110100111" when"111110100101",
"111111110101000" when"111110100110",
"111111110101001" when"111110100111",
"111111110101010" when"111110101000",
"111111110101011" when"111110101001",
"111111110101100" when"111110101010",
"111111110101101" when"111110101011",
"111111110101110" when"111110101100",
"111111110101111" when"111110101101",
"111111110110000" when"111110101110",
"111111110110001" when"111110101111",
"111111110110010" when"111110110000",
"111111110110011" when"111110110001",
"111111110110100" when"111110110010",
"111111110110101" when"111110110011",
"111111110110110" when"111110110100",
"111111110110111" when"111110110101",
"111111110111000" when"111110110110",
"111111110111001" when"111110110111",
"111111110111010" when"111110111000",
"111111110111011" when"111110111001",
"111111110111100" when"111110111010",
"111111110111101" when"111110111011",
"111111110111110" when"111110111100",
"111111110111111" when"111110111101",
"111111111000000" when"111110111110",
"111111111000001" when"111110111111",
"111111111000010" when"111111000000",
"111111111000011" when"111111000001",
"111111111000100" when"111111000010",
"111111111000101" when"111111000011",
"111111111000110" when"111111000100",
"111111111000111" when"111111000101",
"111111111001000" when"111111000110",
"111111111001001" when"111111000111",
"111111111001010" when"111111001000",
"111111111001011" when"111111001001",
"111111111001100" when"111111001010",
"111111111001101" when"111111001011",
"111111111001110" when"111111001100",
"111111111001111" when"111111001101",
"111111111010000" when"111111001110",
"111111111010001" when"111111001111",
"111111111010010" when"111111010000",
"111111111010010" when"111111010001",
"111111111010011" when"111111010010",
"111111111010100" when"111111010011",
"111111111010101" when"111111010100",
"111111111010110" when"111111010101",
"111111111010111" when"111111010110",
"111111111011000" when"111111010111",
"111111111011001" when"111111011000",
"111111111011010" when"111111011001",
"111111111011011" when"111111011010",
"111111111011100" when"111111011011",
"111111111011101" when"111111011100",
"111111111011110" when"111111011101",
"111111111011111" when"111111011110",
"111111111100000" when"111111011111",
"111111111100001" when"111111100000",
"111111111100010" when"111111100001",
"111111111100011" when"111111100010",
"111111111100100" when"111111100011",
"111111111100101" when"111111100100",
"111111111100110" when"111111100101",
"111111111100111" when"111111100110",
"111111111101000" when"111111100111",
"111111111101001" when"111111101000",
"111111111101010" when"111111101001",
"111111111101011" when"111111101010",
"111111111101100" when"111111101011",
"111111111101101" when"111111101100",
"111111111101110" when"111111101101",
"111111111101111" when"111111101110",
"111111111110000" when"111111101111",
"111111111110001" when"111111110000",
"111111111110010" when"111111110001",
"111111111110010" when"111111110010",
"111111111110011" when"111111110011",
"111111111110100" when"111111110100",
"111111111110101" when"111111110101",
"111111111110110" when"111111110110",
"111111111110111" when"111111110111",
"111111111111000" when"111111111000",
"111111111111001" when"111111111001",
"111111111111010" when"111111111010",
"111111111111011" when"111111111011",
"111111111111100" when"111111111100",
"111111111111101" when"111111111101",
"111111111111110" when"111111111110",
"111111111111111" when"111111111111";

end Behavioral;
