 -- 
-- Revision: 1.1: Add several test features
--              Feedback/Fixed output switch (sw[13])
--              3 Fixed outputs(sw[5 downto 3])
--              3 Set points(sw[9 downto 6]) 
--              Inteval switch to swtich between active feedback and slow observation    
--          1.2:
--              Add output threshold. 
--              Remove the inteval switch
--              Fix sensitivity list warnings.
--              2nd: increase the interval time from 10 to 30 cycles.
--          1.3
--              Replace the output switches with treshold switches
--          3.0: 
--              Two channels ad conversion, add an mode switch to distinguish between
--              two photon and florescence. Add another DA output for X. Vaiable
--              "display" is changed to 5 bits to acomodate "2Pho" and "Flor" 
--          5.0:
--              Combine 3.0 and 1.3    
--          5.1:
--              Add the LUT generation function. The lookup table is generated by a
--              block_ram_gene IP
--          6.0:
--              Use the 24bit-12bit division, output log value.  
--          6.1:
--              Use the test switches to configure x output.      
--              Now x_output port will output the RAM value during Lookup table 
--              configuration
--          6.2 Add test configuration.
--              Now during the lookup table generation, a second dac is used to
--              replace the wait state.
--          6.3 LUT gen now goes from 0 to 2*treshold.
--              Now the delay in LUT is performed by repeating DA-AD process.After
--              127 DA-ADs, address increase by '1'.s
--          7.0 Simulation version
--          7.1 Add sync state control of ram reading. The p_in is updated only 
--              during the DAconversion state.
--              Correct the X_outreg assignment problem. 
--          8.0 Implemented new division output argorithm, use two 12-15 bit logs
--              subtraction.
--              Added V_PIDreg to the sensitivity list. 
--          8.1 Now during the LUT gen process, address will hault at 0 for a while
--              to wait for the response of EOM.
--          8.5 Instead of calculating P^2, now log(S) - 2*log(P) is calculated. To
--              do this, log1215 is replaced by log1214, which generates a 14bit 
--              log output. Then, log(P) is left shifted by 1bit, and "11"is added 
--              to log(S).
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity PID is
    Port ( -- system inputs
--           bb0 : out STD_LOGIC_Vector(9 downto 0);
--           bb1 : out STD_LOGIC_Vector(9 downto 0); 
--           input   : out std_logic_vector(11 downto 0);
--           output  : out std_logic_vector(15 downto 0);
           CLK : in STD_LOGIC;
           RST : in STD_LOGIC;
           MODE_SW : in STD_LOGIC;           
           OUT_SW : in STD_LOGIC_VECTOR (2 downto 0);
           TEST_MD : in STD_LOGIC;   
           START : in STD_LOGIC;
           -- IO ports             
           DATA_AD1 : in STD_LOGIC;
           SCLK_AD1 : out STD_LOGIC;
           nCS_AD1 : out STD_LOGIC;
           SCLK_DA3 : out STD_LOGIC;
           nCS_DA3 : out STD_LOGIC;
           nLDAC : out STD_LOGIC;
           DATA_DA3 : out STD_LOGIC;
           SCLK_DA3x : out STD_LOGIC;
           nCS_DA3x : out STD_LOGIC;
           nLDACx : out STD_LOGIC;
           DATA_DA3x : out STD_LOGIC;
           -- 7 segment display ports
           SSEG : out STD_LOGIC_VECTOR (7 downto 0);
           SSAN : out STD_LOGIC_VECTOR (3 downto 0);
           -- Value assignment ports.
           BTN : in STD_LOGIC_VECTOR (1 downto 0);
           INC_SW : in STD_LOGIC_VECTOR (2 downto 0);
           FIX_SW : in STD_LOGIC;
           sw1         : in STD_LOGIC_VECTOR(2 downto 0);
           TRE_SW : in STD_LOGIC;
           LUT_SW : in STD_LOGIC;
           LOG_SW : in STD_LOGIC;
           led  : out STD_LOGIC_VECTOR(15 downto 0)   );
--------------------------------------------------------------------------------
-- Title            : Port Assignments
--
-- Description      : The following signals will be used to drive the  
--                    processes of this VHDL file.
--
--   CLK            : 100MHz on board clock
--
--   RST            : System resets 
--                   
--   MODE_SW        : Control the system state. When '0', system is in test 
--                    running state, when '1', system is in value assignment state
--                   
--   OUT_SW         : Test features. Switch output between input, error, sum 
--                    and pid_out. 
--                   
--   TEST_MD        : Switch between two-photon(1) and florecence(0) imaging
--                   
--   START          : Start pid feedback
--                  
--   BTN            : This is the signal that control the value assignment of 
--                    PID coefficient b0 and b1
--   INC_SW         : This is the vector that corresponds to the three input 
--                    switches that control the increment of the assigned value
--
--   FIX_SW         : This is the switch that controls if the output is a pre-set
--                    value or the PID feedback value.
--
--   sw1            : Test feature. Used for setting different PID set point
--
--   TRE_SW         : This is the switch of turning on/off the output threshold. 
--
--   LUT_SW         : Control the system state. When '0', system is in test 
--                    running state, when '1', system is in Lookup-table-gen
--                    state.
--   LOG_SW         : Test feature. Used to select between log or normal output.
--------------------------------------------------------------------------------        
end PID;

architecture Behavioral of PID is
component assignvalue is
  Port ( 
    RST         : in STD_LOGIC;
    BTN         : in STD_LOGIC_VECTOR (1 downto 0);
    CLK         : in STD_LOGIC;
    en_assign   : in STD_LOGIC;
    SW          : in STD_LOGIC_VECTOR (2 downto 0);
    b1          : out STD_LOGIC_VECTOR (9 downto 0);
    b2          : out STD_LOGIC_VECTOR (9 downto 0);
    out1        : out STD_LOGIC_VECTOR (3 downto 0);
    out2        : out STD_LOGIC_VECTOR (3 downto 0);
    out3        : out STD_LOGIC_VECTOR (3 downto 0));
end component;
component pmodad1 is
  Port    (    
  --General usage
    CLK      : in std_logic;         
    RST      : in std_logic;
     
  --Pmod interface signals
    SDATA    : in std_logic;
    SCLK     : out std_logic;
    nCS      : out std_logic;
        
    --User interface signals
    DATA     : out std_logic_vector(11 downto 0);
    START    : in std_logic; 
    DONE     : out std_logic
            );
end component;
component pmodda3 is
  Port    (    
  --General usage
    CLK      : in std_logic;         
    RST      : in std_logic;
     
  --Pmod interface signals
    DATA     : in std_logic_vector(15 downto 0);
    SCLK     : out std_logic;
    nCS      : out std_logic;
    nLDAC    : out std_logic;
  
  --User interface signals
    INDATA   : out std_logic; 
    START    : in std_logic; 
    start_ad1: in std_logic; 
    DONE     : out std_logic
            );
end component;     

component sseg_display is
    Port ( 
    CLK      : in STD_LOGIC;
    RST      : in STD_LOGIC;
    display1 : in STD_LOGIC_VECTOR (4 downto 0);
    display2 : in STD_LOGIC_VECTOR (4 downto 0);
    display3 : in STD_LOGIC_VECTOR (4 downto 0);
    display4 : in STD_LOGIC_VECTOR (4 downto 0);
    SSEG_CA  : out STD_LOGIC_VECTOR(7 downto 0);
    SSEG_AN  : out STD_LOGIC_VECTOR(3 downto 0));
end component;

component Calculation is
    Port ( DATA_IN  : in STD_LOGIC_VECTOR (11 downto 0);
    P_IN        : in STD_LOGIC_VECTOR (11 downto 0);
    DATA_OUT    : out STD_LOGIC_VECTOR (15 downto 0);
    X_OUT       : out STD_LOGIC_VECTOR (15 downto 0);
    RST         : in STD_LOGIC;
    CLK         : in STD_LOGIC;
    en_reg      : in STD_LOGIC;
    en_cal      : in STD_LOGIC;
    b0          : in STD_LOGIC_VECTOR (9 downto 0);
    b1          : in STD_LOGIC_VECTOR (9 downto 0);
    OUT_SW      : in STD_LOGIC_VECTOR (2 downto 0);
    TEST_MD     : in STD_LOGIC;
    FIX_SW      : in STD_LOGIC;
    sw1         : in STD_LOGIC_VECTOR(2 downto 0);
    TRE_SW      : in STD_LOGIC;
    LOG_SW      : in STD_LOGIC;
    DONE        : out STD_LOGIC);
end component;

component response is
    Port ( CLK : in STD_LOGIC;
           start_rd : in STD_LOGIC;
           done_rd : out STD_LOGIC;
           interval : in STD_LOGIC_VECTOR (23 downto 0));
end component;

COMPONENT power_lut
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(11 DOWNTO 0)
  );
END COMPONENT;

-- A total 4 state are used to control the system       
type states is (Idle,   
                ValueAssign,                
                ADConversion, 
                DataCalculation,
                DAConversion,
                Ready,
                LUTDA,
                LUTAD);                  
signal current_state: states;
signal next_state   : states;

-- start_ad1 signal triggers the AD conversion
-- done_ad1 signal goes high when AD conversion is done and input data vector
-- updated. When a new round of conversion starts, it remains low.
signal start_ad1    : std_logic;
signal done_ad1     : std_logic;
signal start_da3    : std_logic;
signal done_da3     : std_logic;
signal done_da3x    : std_logic;
signal done_cal     : std_logic;
-- control signal for LUT generation
signal en_lut       : std_logic;
-- control signals for value assignment
signal en_assign    : std_logic;
-- control signals for calculation
signal en_reg       : std_logic;
signal en_cal       : std_logic;
-- control signals for ready_wait
signal start_rd     : std_logic;
signal done_rd      : std_logic;
--  registers of value assignment
signal counter1     : STD_LOGIC_VECTOR (3 downto 0);
signal counter2     : STD_LOGIC_VECTOR (3 downto 0);
signal counter3     : STD_LOGIC_VECTOR (3 downto 0);
-- register of 7 segment display
signal display1     : STD_LOGIC_VECTOR (4 downto 0);
signal display2     : STD_LOGIC_VECTOR (4 downto 0);
signal display3     : STD_LOGIC_VECTOR (4 downto 0);
signal display4     : STD_LOGIC_VECTOR (4 downto 0);
-- register of calculation
signal input_data   : std_logic_vector(11 downto 0);
signal p_data       : std_logic_vector(11 downto 0);
signal output_data  : std_logic_vector(15 downto 0);
--signal data_reg     : STD_LOGIC_VECTOR(15 downto 0);
signal dac_data     : std_logic_vector(15 downto 0);
signal x_data       : std_logic_vector(15 downto 0);
signal xdac_data    : std_logic_vector(15 downto 0);
-- PID parameters
signal b0           : STD_LOGIC_VECTOR (9 downto 0);
signal b1           : STD_LOGIC_VECTOR (9 downto 0);
constant interval     : STD_LOGIC_VECTOR (23 downto 0):=x"0000ef";

-- LUT variables
signal address      : STD_LOGIC_VECTOR (15 downto 0):=x"0000";
signal address_s    : STD_LOGIC_VECTOR (14 downto 0):="000000000000000";
--signal lut_counter : STD_LOGIC_VECTOR (31 downto 0):=x"00000001";
signal lut_counter  : STD_LOGIC_VECTOR (6 downto 0):="0000000";
signal zero_pause   : STD_LOGIC;
-- address value of the LUT
signal en_ram       : STD_LOGIC;
-- enable signal of ram
signal en_write     : STD_LOGIC_VECTOR (0 downto 0);
-- enable signal of writing
signal ramin        : STD_LOGIC_VECTOR (11 downto 0);
-- input(recording) signal of ram
signal ramout       : STD_LOGIC_VECTOR (11 downto 0);
-- readout signal of ram

begin

--bb0 <= done_ad1&b0(8 downto 0);
--bb1 <= b1;
--input <= lut_counter&"00000";
--output <= address_s&"0";

-----------------------------------------------------------------------------------
--
-- Title      : Entity Call
--
-- Description: This is the process where the AD converter an DA converter process 
--              are called.
--    
----------------------------------------------------------------------------------- 
    sv: assignvalue port map(        
        RST,
        BTN,
        CLK,
        en_assign,
        INC_SW,
        b0,
        b1,
        counter1,
        counter2,
        counter3);
                   
    adc: pmodad1 port map(   
            CLK,   
            RST,
            DATA_AD1,
            SCLK_AD1,
            nCS_AD1,
            input_data,
            start_ad1,
            done_ad1
                );
                
    cal: Calculation port map(
        input_data,
        p_data,
        output_data,
        x_data,
        RST,
        CLK,
        en_reg,
        en_cal,
        b0,
        b1,
        OUT_SW,
        TEST_MD,
        FIX_SW,
        sw1,        
        TRE_SW,
        LOG_SW,
        done_cal
            );
    dac: pmodda3 port map(
        CLK,         
        RST,
        dac_data,
        SCLK_DA3,
        nCS_DA3,
        nLDAC,
        DATA_DA3, 
        start_da3, 
        start_ad1,
        done_da3
            );

    dacx: pmodda3 port map(
        CLK,         
        RST,
        xdac_data,
        SCLK_DA3x,
        nCS_DA3x,
        nLDACx,
        DATA_DA3x, 
        start_da3, 
        start_ad1,
        done_da3x
            ); 

    sevenseg: sseg_display port map (
        CLK,
        RST,
        display1,
        display2,
        display3,
        display4,
        SSEG,
        SSAN);
    
    wait_response: response port map(
        CLK,
        start_rd,
        done_rd,
        interval);
        
    ram_wr : power_lut PORT MAP (
        clk,
        en_ram,
        en_write,
        address,
        ramin,
        ramout);    
-----------------------------------------------------------------------------------
--
-- Title      : Display Choice
--
-- Description: This is the process were the four digits of the 7 segment dispaly 
--              is assigned. When the system is in the value assignment state, the
--              assigned value and action will show on scree while in the others 
--              states, the display will just show "test".
--
----------------------------------------------------------------------------------- 
display_assignment: process(RST, CLK, en_assign,BTN,START,TEST_MD)
    begin
       if (RST = '1') then
           display1 <= "11111";
           display2 <= "11111";
           display3 <= "11111";
           display4 <= "11111";
       elsif en_assign ='1' then 
       -- when system is in value_assign state
           if BTN(0) = '1' then
           -- when button0 is pressed, counter value is assigned to b0
           display1 <= "01110";
           display2 <= "00000";
           display3 <= "01010";
           display4 <= "11111"; 
           elsif BTN(1) = '1' then
           -- when button0 is pressed, counter value is assigned to b0
           display1 <= "01110";
           display2 <= "00001";
           display3 <= "01010";
           display4 <= "11111";
           else 
           -- when no button is pressed, display the counter value
           display1 <= '0'&counter1;
           display2 <= '0'&counter2;
           display3 <= '0'&counter3;
           display4 <= "11111";
           end if;              
       elsif START = '0' then 
       -- if START switch is low, display "test" to indicate ready
           display1 <= "01100";
           display2 <= "00101";
           display3 <= "01011";
           display4 <= "01100";
       elsif TEST_MD = '0' then
       -- in the florescence state
           display1 <= "10101";
           display2 <= "10011";
           display3 <= "10010";
           display4 <= "10000"; 
       else 
       -- in the two-photon state
           display1 <= "10011";
           display2 <= "10001";
           display3 <= "10100";
           display4 <= "00010";                
       end if;
   end process;  
                
---------------------------------------------------------------------------------
--
-- Title      : Finite State Machine
--
-- Description: A total 9 states are use to control the input/output process.
--              The first state is the Idle state in which the system waits 
--              for the "START" command.
--
--              The second state is the ADConversion state where the pmod ad1
--              takes in analog data and transfer it to digital form. The state
--              is triggerd by the rising edge of signal "start_ad1". At the 
--              end of the state, register "input_data" will be updated and the 
--              signal "done_ad1" will rise.
--
--              The third state is the DataCalculation state. Here no calculation
--              is performed. Instead, "input_data" is right shfited by 4 bits to
--              fit the MSB of the "output_data".
--
--              The fourth state is the DAConversion state in which the data stored
--              in "output_data" is converted. The state is triggerd by the rising
--              edge of "start_da3". "done_da3" will rise when the process is done.
--              The fifth state is ValueAssign state in which the PID coefficient 
--              b0 and b1 is assigned.
--
--              The sixth state is Ready in which is system wait the controlled 
--              to response to the last PID output value.
--
--              The seventh state LUTDA is the DAC process of LUT-generation.
--
--              The eighth state LUTWA is the wait process of LUT-generation.
--
--              The ninth state LUTAD is the ADC process of LUT-generation.
--
-- Notes:       The whole process costs 1700 ns.
--
----------------------------------------------------------------------------------- 
-----------------------------------------------------------------------------------
--
-- Title      : SYNC_PROC
--
-- Description: This is the process were the states are changed synchronously. At 
--              reset the current state becomes Idle state.
--    
-----------------------------------------------------------------------------------            
SYNC_PROC: process (CLK,RST)
   begin
      if (rising_edge(CLK)) then
         if (RST = '1') then
            current_state <= Idle;
         else
            current_state <= next_state;
         end if;        
      end if;
   end process;
    
-----------------------------------------------------------------------------------
--
-- Title      : OUTPUT_DECODE
--
-- Description: This is the process were the output signals are generated
--              unsynchronously based on the state only (Moore State Machine).
--              "en_reg" signal is to enable the update of PID registers, which 
--              should occur before the PID process and only once. So the signal
--              is high in the ADConversion state.
-----------------------------------------------------------------------------------        
OUTPUT_DECODE: process (current_state)
   begin
      if current_state = Idle then
            en_assign <= '0';
            start_ad1 <='0';
            en_cal <= '0';
            en_reg <= '0';
            start_da3 <='0';
            start_rd <= '0';
            en_ram <= '0';            
--            led <= "100000";
        elsif current_state = ValueAssign then
            en_assign <= '1';
            start_ad1 <='0';
            en_cal <= '0';
            en_reg <= '0';
            start_da3 <='0';
            start_rd <= '0';
            en_ram <= '0';            
--            led <= "000001";     
        elsif current_state = ADConversion then
            en_assign <= '0';
            start_ad1 <='1';
            en_cal <= '0';
            en_reg <= '1';
            start_da3 <='0';
            start_rd <= '0';
            en_ram <= '0';
--            led <= "010000";
        elsif current_state = DataCalculation then
            en_assign <= '0';
            start_ad1 <='0';
            en_cal <= '1';
            en_reg <= '0';
            start_da3 <='0';
            start_rd <= '0';
            en_ram <= '0';
--            led <= "001000";            
         elsif current_state = DAConversion then
            en_assign <= '0';
            start_ad1 <='0';
            en_cal <= '0';
            en_reg <= '0';
            start_da3 <='1';
            start_rd <= '0' ;
            en_ram <= '1';
--            led <= "000100";
        elsif current_state = Ready then
            en_assign <= '0';
            start_ad1 <='0';
            en_cal <= '0';
            en_reg <= '0';
            start_da3 <='0';  
            start_rd <= '1'; 
            en_ram <= '0';
--            led <= "000010";           
        elsif current_state = LUTDA then
            en_assign <= '0';
            start_ad1 <='0';
            en_cal <= '0';
            en_reg <= '0';
            start_da3 <='1';
            start_rd <= '0';
            en_ram <= '1';
--            led <= "000011";          
        elsif current_state = LUTAD then        
            en_assign <= '0';
            start_ad1 <='1';
            en_cal <= '0';
            en_reg <= '0';
            start_da3 <='0';
            start_rd <= '0';
            en_ram <= '1';
--            led <= "001100";                                                              
        end if;
    end process;    

-----------------------------------------------------------------------------------
--
-- Title      : LUT Calibration
--
-- Description: This is the process where the Power--Output voltage relation is 
--              calibrated.
-----------------------------------------------------------------------------------   
-----------------------------------------------------------------------------------
--
-- Title      : LUT-GEN Work Flow
--
-- Description: This is the workflow of lookup table. 
--              When RST is released, en_ram is high and the ram is in IDLE state. 
--              
--              When LUT_SW is high, system enters LUT-generation state from IDLE.
--              The first state is LUT DAC where the DAConverter output the current
--              address. At falling edge of done_da3, address will increase by 1.
--
--              Then comes the LUT wait state in which the program pause for a
--              period of time and wait for the system to respond to the output
--              Value.
--              
--              Finally, the LUT ADC state initiate the DA Conversion, en_write is
--              1 at rising edge of done_ad1 and input_data is written into the ram.           
----------------------------------------------------------------------------------- 
    LUT_enable: process(RST, CLK, LUT_SW)
    begin
        if RST = '1' then
            en_lut <= '0';
        elsif rising_edge(CLK) then
            en_lut <= LUT_SW;
        end if;
    end process;
    LUT_cyc: process(RST, done_da3, en_lut)
    begin
        if RST = '1' then
            lut_counter <= "0000000";
        elsif en_lut = '1' then
            if rising_edge(done_da3) then
                lut_counter <= lut_counter + '1';
            end if;
        else lut_counter <= "0000000";
        end if;
    end process;

    counter_incre: process(en_lut, RST, done_ad1, lut_counter)
    begin
        if RST = '1' then
            address_s <= "000000000000000";
            zero_pause <= '0';
        elsif en_lut = '1' then            
            if lut_counter = "1111111" then
                if falling_edge(done_ad1) then
                    address_s <= address_s + '1';
                    if address_s = "000000000000000" then
                        zero_pause <= not zero_pause;
                    end if;
                end if;
            end if;
        end if;
    end process;
    
    address_assign: process(RST, en_lut, address_s, zero_pause, start_ad1,output_data)
    begin
        if RST = '1' then
            address <= x"0000";
        elsif en_lut = '1' then
            if zero_pause = '0' then
                address <= '0'&address_s;
            else address <= x"0000";
            end if;
        elsif rising_edge(start_ad1) then
        -- for reading the Lookup table data
            address <= output_data;            
        end if;        
    end process;
    
    with en_lut select dac_data <=
        output_data when '0',
        address      when '1';

    with en_lut select xdac_data <=
        x_data when '0',
        ramout&"0000"   when '1';
                
    led<=xdac_data;

            
    write_ram: process(en_lut, done_ad1)
    begin
        if en_lut = '1' then
            en_write(0) <= done_ad1;
        else en_write <= "0";
        end if;
    end process;
    
    power_assign: process(en_lut,done_ad1)
    begin
        if en_lut = '1' then
            if rising_edge(done_ad1) then
                ramin <= input_data;
            end if;
        end if;
    end process;
    
    power_lookup: process(en_lut, ramout)
    begin
        if en_lut = '0' then
            p_data <= ramout;
        end if;
    end process;                

        
----------------------------------------------------------------------------------
--
-- Title      : NEXT_STATE_DECODE
--
-- Description: This is the process were the next state logic is generated 
--              depending on the current state and the input signals.
--    
-----------------------------------------------------------------------------------    
    NEXT_STATE_DECODE: process (current_state, START, MODE_SW, done_ad1, done_cal, done_da3, done_rd, en_lut)
    begin      
      next_state <= current_state;  -- default is to stay in current state     
      case (current_state) is
         when Idle =>
            if START = '1' then
                next_state <= ADConversion;
            elsif MODE_SW = '1' then
                next_state <= ValueAssign;
            elsif en_lut = '1' then
                next_state <= LUTDA;
            end if;
         when ValueAssign =>
            if MODE_SW = '0' then
                next_state <= Idle;
            end if;                                 
         when ADConversion =>
            if rising_edge(done_ad1) then
               next_state <= DataCalculation;
            end if;
         when DataCalculation =>
            if rising_edge(done_cal) then
                next_state <= DAConversion;
            end if;
         when DAConversion =>
            if rising_edge(done_da3) then
                next_state <= Ready;
            end if;
         when Ready =>
            if rising_edge(done_rd) then
                next_state <= Idle;
            end if;         
         when LUTDA =>
            if rising_edge(done_da3) then
                next_state <= LUTAD;
            end if;        
         when LUTAD =>
            if rising_edge(done_ad1) then
                if en_lut = '1' then   
                    next_state <= LUTDA;
                else
                    next_state <= Idle;
                end if;  
            end if;             
         when others =>
            next_state <= Idle;
      end case;      
   end process;

end Behavioral;
